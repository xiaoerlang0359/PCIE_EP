///////////////////////////////////////////////////////
//  Copyright (c) 2011 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /     Vendor      : Xilinx 
// \  \    \/      Version : 10.1
//  \  \           Description : 
//  /  /                      
// /__/   /\       Filename    : BUFG_LB.v
// \  \  /  \ 
//  \__\/\__ \                    
//                                 
//  Generated by :	/home/unified/patrickp/HEAD/env/Databases/CAEInterfaces/LibraryWriters/bin/ltw.pl
//  Revision:		1.0
//    11/15/11 - 634082 - connected ouput.
//    05/22/12 - 661573 - remove 100 ps delay on output.
//  End Revision
///////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

module BUFG_LB (
  CLKOUT,

  CLKIN
);


  output CLKOUT;

  input CLKIN;

  initial begin
  end

  buf B_CLKOUT (CLKOUT, CLKIN);

  specify
    ( CLKIN *> CLKOUT) = (0, 0);

    specparam PATHPULSE$ = 0;
  endspecify
endmodule
