///////////////////////////////////////////////////////
//  Copyright (c) 2011 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /     Vendor      : Xilinx 
// \  \    \/      Version     : 13.3
//  \  \           Description : 
//  /  /                      
// /__/   /\       Filename    : X_PCIE_3_0.v
// \  \  /  \ 
//  \__\/\__ \                    
//                                 
//  Revision:		1.0
//  02/23/11 - Intial Version : 10.1
//  04/13/11 - 605801 - Updated YML
//  04/28/11 - 608328 - Updated YML & initial secureip publish
//  07/20/11 - 617638 - Updated YML (new attributes)
//  07/26/11 - 618494 - Updated YML
//  01/18/13 - 695630 - added drp monitor
///////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

module X_PCIE_3_0 (
  CFGCURRENTSPEED,
  CFGDPASUBSTATECHANGE,
  CFGERRCOROUT,
  CFGERRFATALOUT,
  CFGERRNONFATALOUT,
  CFGEXTFUNCTIONNUMBER,
  CFGEXTREADRECEIVED,
  CFGEXTREGISTERNUMBER,
  CFGEXTWRITEBYTEENABLE,
  CFGEXTWRITEDATA,
  CFGEXTWRITERECEIVED,
  CFGFCCPLD,
  CFGFCCPLH,
  CFGFCNPD,
  CFGFCNPH,
  CFGFCPD,
  CFGFCPH,
  CFGFLRINPROCESS,
  CFGFUNCTIONPOWERSTATE,
  CFGFUNCTIONSTATUS,
  CFGHOTRESETOUT,
  CFGINPUTUPDATEDONE,
  CFGINTERRUPTAOUTPUT,
  CFGINTERRUPTBOUTPUT,
  CFGINTERRUPTCOUTPUT,
  CFGINTERRUPTDOUTPUT,
  CFGINTERRUPTMSIDATA,
  CFGINTERRUPTMSIENABLE,
  CFGINTERRUPTMSIFAIL,
  CFGINTERRUPTMSIMASKUPDATE,
  CFGINTERRUPTMSIMMENABLE,
  CFGINTERRUPTMSISENT,
  CFGINTERRUPTMSIVFENABLE,
  CFGINTERRUPTMSIXENABLE,
  CFGINTERRUPTMSIXFAIL,
  CFGINTERRUPTMSIXMASK,
  CFGINTERRUPTMSIXSENT,
  CFGINTERRUPTMSIXVFENABLE,
  CFGINTERRUPTMSIXVFMASK,
  CFGINTERRUPTSENT,
  CFGLINKPOWERSTATE,
  CFGLOCALERROR,
  CFGLTRENABLE,
  CFGLTSSMSTATE,
  CFGMAXPAYLOAD,
  CFGMAXREADREQ,
  CFGMCUPDATEDONE,
  CFGMGMTREADDATA,
  CFGMGMTREADWRITEDONE,
  CFGMSGRECEIVED,
  CFGMSGRECEIVEDDATA,
  CFGMSGRECEIVEDTYPE,
  CFGMSGTRANSMITDONE,
  CFGNEGOTIATEDWIDTH,
  CFGOBFFENABLE,
  CFGPERFUNCSTATUSDATA,
  CFGPERFUNCTIONUPDATEDONE,
  CFGPHYLINKDOWN,
  CFGPHYLINKSTATUS,
  CFGPLSTATUSCHANGE,
  CFGPOWERSTATECHANGEINTERRUPT,
  CFGRCBSTATUS,
  CFGTPHFUNCTIONNUM,
  CFGTPHREQUESTERENABLE,
  CFGTPHSTMODE,
  CFGTPHSTTADDRESS,
  CFGTPHSTTREADENABLE,
  CFGTPHSTTWRITEBYTEVALID,
  CFGTPHSTTWRITEDATA,
  CFGTPHSTTWRITEENABLE,
  CFGVFFLRINPROCESS,
  CFGVFPOWERSTATE,
  CFGVFSTATUS,
  CFGVFTPHREQUESTERENABLE,
  CFGVFTPHSTMODE,
  DBGDATAOUT,
  DRPDO,
  DRPRDY,
  MAXISCQTDATA,
  MAXISCQTKEEP,
  MAXISCQTLAST,
  MAXISCQTUSER,
  MAXISCQTVALID,
  MAXISRCTDATA,
  MAXISRCTKEEP,
  MAXISRCTLAST,
  MAXISRCTUSER,
  MAXISRCTVALID,
  MICOMPLETIONRAMREADADDRESSAL,
  MICOMPLETIONRAMREADADDRESSAU,
  MICOMPLETIONRAMREADADDRESSBL,
  MICOMPLETIONRAMREADADDRESSBU,
  MICOMPLETIONRAMREADENABLEL,
  MICOMPLETIONRAMREADENABLEU,
  MICOMPLETIONRAMWRITEADDRESSAL,
  MICOMPLETIONRAMWRITEADDRESSAU,
  MICOMPLETIONRAMWRITEADDRESSBL,
  MICOMPLETIONRAMWRITEADDRESSBU,
  MICOMPLETIONRAMWRITEDATAL,
  MICOMPLETIONRAMWRITEDATAU,
  MICOMPLETIONRAMWRITEENABLEL,
  MICOMPLETIONRAMWRITEENABLEU,
  MIREPLAYRAMADDRESS,
  MIREPLAYRAMREADENABLE,
  MIREPLAYRAMWRITEDATA,
  MIREPLAYRAMWRITEENABLE,
  MIREQUESTRAMREADADDRESSA,
  MIREQUESTRAMREADADDRESSB,
  MIREQUESTRAMREADENABLE,
  MIREQUESTRAMWRITEADDRESSA,
  MIREQUESTRAMWRITEADDRESSB,
  MIREQUESTRAMWRITEDATA,
  MIREQUESTRAMWRITEENABLE,
  PCIECQNPREQCOUNT,
  PCIERQSEQNUM,
  PCIERQSEQNUMVLD,
  PCIERQTAG,
  PCIERQTAGAV,
  PCIERQTAGVLD,
  PCIETFCNPDAV,
  PCIETFCNPHAV,
  PIPERX0EQCONTROL,
  PIPERX0EQLPLFFS,
  PIPERX0EQLPTXPRESET,
  PIPERX0EQPRESET,
  PIPERX0POLARITY,
  PIPERX1EQCONTROL,
  PIPERX1EQLPLFFS,
  PIPERX1EQLPTXPRESET,
  PIPERX1EQPRESET,
  PIPERX1POLARITY,
  PIPERX2EQCONTROL,
  PIPERX2EQLPLFFS,
  PIPERX2EQLPTXPRESET,
  PIPERX2EQPRESET,
  PIPERX2POLARITY,
  PIPERX3EQCONTROL,
  PIPERX3EQLPLFFS,
  PIPERX3EQLPTXPRESET,
  PIPERX3EQPRESET,
  PIPERX3POLARITY,
  PIPERX4EQCONTROL,
  PIPERX4EQLPLFFS,
  PIPERX4EQLPTXPRESET,
  PIPERX4EQPRESET,
  PIPERX4POLARITY,
  PIPERX5EQCONTROL,
  PIPERX5EQLPLFFS,
  PIPERX5EQLPTXPRESET,
  PIPERX5EQPRESET,
  PIPERX5POLARITY,
  PIPERX6EQCONTROL,
  PIPERX6EQLPLFFS,
  PIPERX6EQLPTXPRESET,
  PIPERX6EQPRESET,
  PIPERX6POLARITY,
  PIPERX7EQCONTROL,
  PIPERX7EQLPLFFS,
  PIPERX7EQLPTXPRESET,
  PIPERX7EQPRESET,
  PIPERX7POLARITY,
  PIPETX0CHARISK,
  PIPETX0COMPLIANCE,
  PIPETX0DATA,
  PIPETX0DATAVALID,
  PIPETX0ELECIDLE,
  PIPETX0EQCONTROL,
  PIPETX0EQDEEMPH,
  PIPETX0EQPRESET,
  PIPETX0POWERDOWN,
  PIPETX0STARTBLOCK,
  PIPETX0SYNCHEADER,
  PIPETX1CHARISK,
  PIPETX1COMPLIANCE,
  PIPETX1DATA,
  PIPETX1DATAVALID,
  PIPETX1ELECIDLE,
  PIPETX1EQCONTROL,
  PIPETX1EQDEEMPH,
  PIPETX1EQPRESET,
  PIPETX1POWERDOWN,
  PIPETX1STARTBLOCK,
  PIPETX1SYNCHEADER,
  PIPETX2CHARISK,
  PIPETX2COMPLIANCE,
  PIPETX2DATA,
  PIPETX2DATAVALID,
  PIPETX2ELECIDLE,
  PIPETX2EQCONTROL,
  PIPETX2EQDEEMPH,
  PIPETX2EQPRESET,
  PIPETX2POWERDOWN,
  PIPETX2STARTBLOCK,
  PIPETX2SYNCHEADER,
  PIPETX3CHARISK,
  PIPETX3COMPLIANCE,
  PIPETX3DATA,
  PIPETX3DATAVALID,
  PIPETX3ELECIDLE,
  PIPETX3EQCONTROL,
  PIPETX3EQDEEMPH,
  PIPETX3EQPRESET,
  PIPETX3POWERDOWN,
  PIPETX3STARTBLOCK,
  PIPETX3SYNCHEADER,
  PIPETX4CHARISK,
  PIPETX4COMPLIANCE,
  PIPETX4DATA,
  PIPETX4DATAVALID,
  PIPETX4ELECIDLE,
  PIPETX4EQCONTROL,
  PIPETX4EQDEEMPH,
  PIPETX4EQPRESET,
  PIPETX4POWERDOWN,
  PIPETX4STARTBLOCK,
  PIPETX4SYNCHEADER,
  PIPETX5CHARISK,
  PIPETX5COMPLIANCE,
  PIPETX5DATA,
  PIPETX5DATAVALID,
  PIPETX5ELECIDLE,
  PIPETX5EQCONTROL,
  PIPETX5EQDEEMPH,
  PIPETX5EQPRESET,
  PIPETX5POWERDOWN,
  PIPETX5STARTBLOCK,
  PIPETX5SYNCHEADER,
  PIPETX6CHARISK,
  PIPETX6COMPLIANCE,
  PIPETX6DATA,
  PIPETX6DATAVALID,
  PIPETX6ELECIDLE,
  PIPETX6EQCONTROL,
  PIPETX6EQDEEMPH,
  PIPETX6EQPRESET,
  PIPETX6POWERDOWN,
  PIPETX6STARTBLOCK,
  PIPETX6SYNCHEADER,
  PIPETX7CHARISK,
  PIPETX7COMPLIANCE,
  PIPETX7DATA,
  PIPETX7DATAVALID,
  PIPETX7ELECIDLE,
  PIPETX7EQCONTROL,
  PIPETX7EQDEEMPH,
  PIPETX7EQPRESET,
  PIPETX7POWERDOWN,
  PIPETX7STARTBLOCK,
  PIPETX7SYNCHEADER,
  PIPETXDEEMPH,
  PIPETXMARGIN,
  PIPETXRATE,
  PIPETXRCVRDET,
  PIPETXRESET,
  PIPETXSWING,
  PLEQINPROGRESS,
  PLEQPHASE,
  PLGEN3PCSRXSLIDE,
  SAXISCCTREADY,
  SAXISRQTREADY,

  CFGCONFIGSPACEENABLE,
  CFGDEVID,
  CFGDSBUSNUMBER,
  CFGDSDEVICENUMBER,
  CFGDSFUNCTIONNUMBER,
  CFGDSN,
  CFGDSPORTNUMBER,
  CFGERRCORIN,
  CFGERRUNCORIN,
  CFGEXTREADDATA,
  CFGEXTREADDATAVALID,
  CFGFCSEL,
  CFGFLRDONE,
  CFGHOTRESETIN,
  CFGINPUTUPDATEREQUEST,
  CFGINTERRUPTINT,
  CFGINTERRUPTMSIATTR,
  CFGINTERRUPTMSIFUNCTIONNUMBER,
  CFGINTERRUPTMSIINT,
  CFGINTERRUPTMSIPENDINGSTATUS,
  CFGINTERRUPTMSISELECT,
  CFGINTERRUPTMSITPHPRESENT,
  CFGINTERRUPTMSITPHSTTAG,
  CFGINTERRUPTMSITPHTYPE,
  CFGINTERRUPTMSIXADDRESS,
  CFGINTERRUPTMSIXDATA,
  CFGINTERRUPTMSIXINT,
  CFGINTERRUPTPENDING,
  CFGLINKTRAININGENABLE,
  CFGMCUPDATEREQUEST,
  CFGMGMTADDR,
  CFGMGMTBYTEENABLE,
  CFGMGMTREAD,
  CFGMGMTTYPE1CFGREGACCESS,
  CFGMGMTWRITE,
  CFGMGMTWRITEDATA,
  CFGMSGTRANSMIT,
  CFGMSGTRANSMITDATA,
  CFGMSGTRANSMITTYPE,
  CFGPERFUNCSTATUSCONTROL,
  CFGPERFUNCTIONNUMBER,
  CFGPERFUNCTIONOUTPUTREQUEST,
  CFGPOWERSTATECHANGEACK,
  CFGREQPMTRANSITIONL23READY,
  CFGREVID,
  CFGSUBSYSID,
  CFGSUBSYSVENDID,
  CFGTPHSTTREADDATA,
  CFGTPHSTTREADDATAVALID,
  CFGVENDID,
  CFGVFFLRDONE,
  CORECLK,
  CORECLKMICOMPLETIONRAML,
  CORECLKMICOMPLETIONRAMU,
  CORECLKMIREPLAYRAM,
  CORECLKMIREQUESTRAM,
  DRPADDR,
  DRPCLK,
  DRPDI,
  DRPEN,
  DRPWE,
  MAXISCQTREADY,
  MAXISRCTREADY,
  MGMTRESETN,
  MGMTSTICKYRESETN,
  MICOMPLETIONRAMREADDATA,
  MIREPLAYRAMREADDATA,
  MIREQUESTRAMREADDATA,
  PCIECQNPREQ,
  PIPECLK,
  PIPEEQFS,
  PIPEEQLF,
  PIPERESETN,
  PIPERX0CHARISK,
  PIPERX0DATA,
  PIPERX0DATAVALID,
  PIPERX0ELECIDLE,
  PIPERX0EQDONE,
  PIPERX0EQLPADAPTDONE,
  PIPERX0EQLPLFFSSEL,
  PIPERX0EQLPNEWTXCOEFFORPRESET,
  PIPERX0PHYSTATUS,
  PIPERX0STARTBLOCK,
  PIPERX0STATUS,
  PIPERX0SYNCHEADER,
  PIPERX0VALID,
  PIPERX1CHARISK,
  PIPERX1DATA,
  PIPERX1DATAVALID,
  PIPERX1ELECIDLE,
  PIPERX1EQDONE,
  PIPERX1EQLPADAPTDONE,
  PIPERX1EQLPLFFSSEL,
  PIPERX1EQLPNEWTXCOEFFORPRESET,
  PIPERX1PHYSTATUS,
  PIPERX1STARTBLOCK,
  PIPERX1STATUS,
  PIPERX1SYNCHEADER,
  PIPERX1VALID,
  PIPERX2CHARISK,
  PIPERX2DATA,
  PIPERX2DATAVALID,
  PIPERX2ELECIDLE,
  PIPERX2EQDONE,
  PIPERX2EQLPADAPTDONE,
  PIPERX2EQLPLFFSSEL,
  PIPERX2EQLPNEWTXCOEFFORPRESET,
  PIPERX2PHYSTATUS,
  PIPERX2STARTBLOCK,
  PIPERX2STATUS,
  PIPERX2SYNCHEADER,
  PIPERX2VALID,
  PIPERX3CHARISK,
  PIPERX3DATA,
  PIPERX3DATAVALID,
  PIPERX3ELECIDLE,
  PIPERX3EQDONE,
  PIPERX3EQLPADAPTDONE,
  PIPERX3EQLPLFFSSEL,
  PIPERX3EQLPNEWTXCOEFFORPRESET,
  PIPERX3PHYSTATUS,
  PIPERX3STARTBLOCK,
  PIPERX3STATUS,
  PIPERX3SYNCHEADER,
  PIPERX3VALID,
  PIPERX4CHARISK,
  PIPERX4DATA,
  PIPERX4DATAVALID,
  PIPERX4ELECIDLE,
  PIPERX4EQDONE,
  PIPERX4EQLPADAPTDONE,
  PIPERX4EQLPLFFSSEL,
  PIPERX4EQLPNEWTXCOEFFORPRESET,
  PIPERX4PHYSTATUS,
  PIPERX4STARTBLOCK,
  PIPERX4STATUS,
  PIPERX4SYNCHEADER,
  PIPERX4VALID,
  PIPERX5CHARISK,
  PIPERX5DATA,
  PIPERX5DATAVALID,
  PIPERX5ELECIDLE,
  PIPERX5EQDONE,
  PIPERX5EQLPADAPTDONE,
  PIPERX5EQLPLFFSSEL,
  PIPERX5EQLPNEWTXCOEFFORPRESET,
  PIPERX5PHYSTATUS,
  PIPERX5STARTBLOCK,
  PIPERX5STATUS,
  PIPERX5SYNCHEADER,
  PIPERX5VALID,
  PIPERX6CHARISK,
  PIPERX6DATA,
  PIPERX6DATAVALID,
  PIPERX6ELECIDLE,
  PIPERX6EQDONE,
  PIPERX6EQLPADAPTDONE,
  PIPERX6EQLPLFFSSEL,
  PIPERX6EQLPNEWTXCOEFFORPRESET,
  PIPERX6PHYSTATUS,
  PIPERX6STARTBLOCK,
  PIPERX6STATUS,
  PIPERX6SYNCHEADER,
  PIPERX6VALID,
  PIPERX7CHARISK,
  PIPERX7DATA,
  PIPERX7DATAVALID,
  PIPERX7ELECIDLE,
  PIPERX7EQDONE,
  PIPERX7EQLPADAPTDONE,
  PIPERX7EQLPLFFSSEL,
  PIPERX7EQLPNEWTXCOEFFORPRESET,
  PIPERX7PHYSTATUS,
  PIPERX7STARTBLOCK,
  PIPERX7STATUS,
  PIPERX7SYNCHEADER,
  PIPERX7VALID,
  PIPETX0EQCOEFF,
  PIPETX0EQDONE,
  PIPETX1EQCOEFF,
  PIPETX1EQDONE,
  PIPETX2EQCOEFF,
  PIPETX2EQDONE,
  PIPETX3EQCOEFF,
  PIPETX3EQDONE,
  PIPETX4EQCOEFF,
  PIPETX4EQDONE,
  PIPETX5EQCOEFF,
  PIPETX5EQDONE,
  PIPETX6EQCOEFF,
  PIPETX6EQDONE,
  PIPETX7EQCOEFF,
  PIPETX7EQDONE,
  PLDISABLESCRAMBLER,
  PLEQRESETEIEOSCOUNT,
  PLGEN3PCSDISABLE,
  PLGEN3PCSRXSYNCDONE,
  RECCLK,
  RESETN,
  SAXISCCTDATA,
  SAXISCCTKEEP,
  SAXISCCTLAST,
  SAXISCCTUSER,
  SAXISCCTVALID,
  SAXISRQTDATA,
  SAXISRQTKEEP,
  SAXISRQTLAST,
  SAXISRQTUSER,
  SAXISRQTVALID,
  USERCLK
);

  parameter LOC = "UNPLACED";
  parameter ARI_CAP_ENABLE = "FALSE";
  parameter AXISTEN_IF_CC_ALIGNMENT_MODE = "FALSE";
  parameter AXISTEN_IF_CC_PARITY_CHK = "TRUE";
  parameter AXISTEN_IF_CQ_ALIGNMENT_MODE = "FALSE";
  parameter AXISTEN_IF_ENABLE_CLIENT_TAG = "FALSE";
  parameter [17:0] AXISTEN_IF_ENABLE_MSG_ROUTE = 18'h00000;
  parameter AXISTEN_IF_ENABLE_RX_MSG_INTFC = "FALSE";
  parameter AXISTEN_IF_RC_ALIGNMENT_MODE = "FALSE";
  parameter AXISTEN_IF_RC_STRADDLE = "FALSE";
  parameter AXISTEN_IF_RQ_ALIGNMENT_MODE = "FALSE";
  parameter AXISTEN_IF_RQ_PARITY_CHK = "TRUE";
  parameter [1:0] AXISTEN_IF_WIDTH = 2'h2;
  parameter CRM_CORE_CLK_FREQ_500 = "TRUE";
  parameter [1:0] CRM_USER_CLK_FREQ = 2'h2;
  parameter [7:0] DNSTREAM_LINK_NUM = 8'h00;
  parameter [1:0] GEN3_PCS_AUTO_REALIGN = 2'h1;
  parameter GEN3_PCS_RX_ELECIDLE_INTERNAL = "TRUE";
  parameter [8:0] LL_ACK_TIMEOUT = 9'h000;
  parameter LL_ACK_TIMEOUT_EN = "FALSE";
  parameter integer LL_ACK_TIMEOUT_FUNC = 0;
  parameter [15:0] LL_CPL_FC_UPDATE_TIMER = 16'h0000;
  parameter LL_CPL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
  parameter [15:0] LL_FC_UPDATE_TIMER = 16'h0000;
  parameter LL_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
  parameter [15:0] LL_NP_FC_UPDATE_TIMER = 16'h0000;
  parameter LL_NP_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
  parameter [15:0] LL_P_FC_UPDATE_TIMER = 16'h0000;
  parameter LL_P_FC_UPDATE_TIMER_OVERRIDE = "FALSE";
  parameter [8:0] LL_REPLAY_TIMEOUT = 9'h000;
  parameter LL_REPLAY_TIMEOUT_EN = "FALSE";
  parameter integer LL_REPLAY_TIMEOUT_FUNC = 0;
  parameter [9:0] LTR_TX_MESSAGE_MINIMUM_INTERVAL = 10'h0FA;
  parameter LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE = "FALSE";
  parameter LTR_TX_MESSAGE_ON_LTR_ENABLE = "FALSE";
  parameter PF0_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
  parameter PF0_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
  parameter [11:0] PF0_AER_CAP_NEXTPTR = 12'h000;
  parameter [11:0] PF0_ARI_CAP_NEXTPTR = 12'h000;
  parameter [7:0] PF0_ARI_CAP_NEXT_FUNC = 8'h00;
  parameter [3:0] PF0_ARI_CAP_VER = 4'h1;
  parameter [4:0] PF0_BAR0_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_BAR0_CONTROL = 3'h4;
  parameter [4:0] PF0_BAR1_APERTURE_SIZE = 5'h00;
  parameter [2:0] PF0_BAR1_CONTROL = 3'h0;
  parameter [4:0] PF0_BAR2_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_BAR2_CONTROL = 3'h4;
  parameter [4:0] PF0_BAR3_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_BAR3_CONTROL = 3'h0;
  parameter [4:0] PF0_BAR4_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_BAR4_CONTROL = 3'h4;
  parameter [4:0] PF0_BAR5_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_BAR5_CONTROL = 3'h0;
  parameter [7:0] PF0_BIST_REGISTER = 8'h00;
  parameter [7:0] PF0_CAPABILITY_POINTER = 8'h50;
  parameter [23:0] PF0_CLASS_CODE = 24'h000000;
  parameter [15:0] PF0_DEVICE_ID = 16'h0000;
  parameter PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT = "TRUE";
  parameter PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
  parameter PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT = "TRUE";
  parameter PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE = "TRUE";
  parameter PF0_DEV_CAP2_LTR_SUPPORT = "TRUE";
  parameter [1:0] PF0_DEV_CAP2_OBFF_SUPPORT = 2'h0;
  parameter PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT = "FALSE";
  parameter integer PF0_DEV_CAP_ENDPOINT_L0S_LATENCY = 0;
  parameter integer PF0_DEV_CAP_ENDPOINT_L1_LATENCY = 0;
  parameter PF0_DEV_CAP_EXT_TAG_SUPPORTED = "TRUE";
  parameter PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE = "TRUE";
  parameter [2:0] PF0_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
  parameter [11:0] PF0_DPA_CAP_NEXTPTR = 12'h000;
  parameter [4:0] PF0_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
  parameter PF0_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
  parameter [7:0] PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
  parameter [3:0] PF0_DPA_CAP_VER = 4'h1;
  parameter [11:0] PF0_DSN_CAP_NEXTPTR = 12'h10C;
  parameter [4:0] PF0_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
  parameter PF0_EXPANSION_ROM_ENABLE = "FALSE";
  parameter [7:0] PF0_INTERRUPT_LINE = 8'h00;
  parameter [2:0] PF0_INTERRUPT_PIN = 3'h1;
  parameter integer PF0_LINK_CAP_ASPM_SUPPORT = 0;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 = 7;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 = 7;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 = 7;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 = 7;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 = 7;
  parameter integer PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 = 7;
  parameter integer PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 = 7;
  parameter PF0_LINK_STATUS_SLOT_CLOCK_CONFIG = "TRUE";
  parameter [9:0] PF0_LTR_CAP_MAX_NOSNOOP_LAT = 10'h000;
  parameter [9:0] PF0_LTR_CAP_MAX_SNOOP_LAT = 10'h000;
  parameter [11:0] PF0_LTR_CAP_NEXTPTR = 12'h000;
  parameter [3:0] PF0_LTR_CAP_VER = 4'h1;
  parameter [7:0] PF0_MSIX_CAP_NEXTPTR = 8'h00;
  parameter integer PF0_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] PF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer PF0_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] PF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] PF0_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer PF0_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] PF0_MSI_CAP_NEXTPTR = 8'h00;
  parameter [11:0] PF0_PB_CAP_NEXTPTR = 12'h000;
  parameter PF0_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
  parameter [3:0] PF0_PB_CAP_VER = 4'h1;
  parameter [7:0] PF0_PM_CAP_ID = 8'h01;
  parameter [7:0] PF0_PM_CAP_NEXTPTR = 8'h00;
  parameter PF0_PM_CAP_PMESUPPORT_D0 = "TRUE";
  parameter PF0_PM_CAP_PMESUPPORT_D1 = "TRUE";
  parameter PF0_PM_CAP_PMESUPPORT_D3HOT = "TRUE";
  parameter PF0_PM_CAP_SUPP_D1_STATE = "TRUE";
  parameter [2:0] PF0_PM_CAP_VER_ID = 3'h3;
  parameter PF0_PM_CSR_NOSOFTRESET = "TRUE";
  parameter PF0_RBAR_CAP_ENABLE = "FALSE";
  parameter [2:0] PF0_RBAR_CAP_INDEX0 = 3'h0;
  parameter [2:0] PF0_RBAR_CAP_INDEX1 = 3'h0;
  parameter [2:0] PF0_RBAR_CAP_INDEX2 = 3'h0;
  parameter [11:0] PF0_RBAR_CAP_NEXTPTR = 12'h000;
  parameter [19:0] PF0_RBAR_CAP_SIZE0 = 20'h00000;
  parameter [19:0] PF0_RBAR_CAP_SIZE1 = 20'h00000;
  parameter [19:0] PF0_RBAR_CAP_SIZE2 = 20'h00000;
  parameter [3:0] PF0_RBAR_CAP_VER = 4'h1;
  parameter [2:0] PF0_RBAR_NUM = 3'h1;
  parameter [7:0] PF0_REVISION_ID = 8'h00;
  parameter [4:0] PF0_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_SRIOV_BAR0_CONTROL = 3'h4;
  parameter [4:0] PF0_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
  parameter [2:0] PF0_SRIOV_BAR1_CONTROL = 3'h0;
  parameter [4:0] PF0_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_SRIOV_BAR2_CONTROL = 3'h4;
  parameter [4:0] PF0_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_SRIOV_BAR3_CONTROL = 3'h0;
  parameter [4:0] PF0_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_SRIOV_BAR4_CONTROL = 3'h4;
  parameter [4:0] PF0_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF0_SRIOV_BAR5_CONTROL = 3'h0;
  parameter [15:0] PF0_SRIOV_CAP_INITIAL_VF = 16'h0000;
  parameter [11:0] PF0_SRIOV_CAP_NEXTPTR = 12'h000;
  parameter [15:0] PF0_SRIOV_CAP_TOTAL_VF = 16'h0000;
  parameter [3:0] PF0_SRIOV_CAP_VER = 4'h1;
  parameter [15:0] PF0_SRIOV_FIRST_VF_OFFSET = 16'h0000;
  parameter [15:0] PF0_SRIOV_FUNC_DEP_LINK = 16'h0000;
  parameter [31:0] PF0_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
  parameter [15:0] PF0_SRIOV_VF_DEVICE_ID = 16'h0000;
  parameter [15:0] PF0_SUBSYSTEM_ID = 16'h0000;
  parameter PF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter PF0_TPHR_CAP_ENABLE = "FALSE";
  parameter PF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] PF0_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] PF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] PF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] PF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] PF0_TPHR_CAP_VER = 4'h1;
  parameter [11:0] PF0_VC_CAP_NEXTPTR = 12'h000;
  parameter [3:0] PF0_VC_CAP_VER = 4'h1;
  parameter PF1_AER_CAP_ECRC_CHECK_CAPABLE = "FALSE";
  parameter PF1_AER_CAP_ECRC_GEN_CAPABLE = "FALSE";
  parameter [11:0] PF1_AER_CAP_NEXTPTR = 12'h000;
  parameter [11:0] PF1_ARI_CAP_NEXTPTR = 12'h000;
  parameter [7:0] PF1_ARI_CAP_NEXT_FUNC = 8'h00;
  parameter [4:0] PF1_BAR0_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_BAR0_CONTROL = 3'h4;
  parameter [4:0] PF1_BAR1_APERTURE_SIZE = 5'h00;
  parameter [2:0] PF1_BAR1_CONTROL = 3'h0;
  parameter [4:0] PF1_BAR2_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_BAR2_CONTROL = 3'h4;
  parameter [4:0] PF1_BAR3_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_BAR3_CONTROL = 3'h0;
  parameter [4:0] PF1_BAR4_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_BAR4_CONTROL = 3'h4;
  parameter [4:0] PF1_BAR5_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_BAR5_CONTROL = 3'h0;
  parameter [7:0] PF1_BIST_REGISTER = 8'h00;
  parameter [7:0] PF1_CAPABILITY_POINTER = 8'h50;
  parameter [23:0] PF1_CLASS_CODE = 24'h000000;
  parameter [15:0] PF1_DEVICE_ID = 16'h0000;
  parameter [2:0] PF1_DEV_CAP_MAX_PAYLOAD_SIZE = 3'h3;
  parameter [11:0] PF1_DPA_CAP_NEXTPTR = 12'h000;
  parameter [4:0] PF1_DPA_CAP_SUB_STATE_CONTROL = 5'h00;
  parameter PF1_DPA_CAP_SUB_STATE_CONTROL_EN = "TRUE";
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 = 8'h00;
  parameter [7:0] PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 = 8'h00;
  parameter [3:0] PF1_DPA_CAP_VER = 4'h1;
  parameter [11:0] PF1_DSN_CAP_NEXTPTR = 12'h10C;
  parameter [4:0] PF1_EXPANSION_ROM_APERTURE_SIZE = 5'h03;
  parameter PF1_EXPANSION_ROM_ENABLE = "FALSE";
  parameter [7:0] PF1_INTERRUPT_LINE = 8'h00;
  parameter [2:0] PF1_INTERRUPT_PIN = 3'h1;
  parameter [7:0] PF1_MSIX_CAP_NEXTPTR = 8'h00;
  parameter integer PF1_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] PF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer PF1_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] PF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] PF1_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer PF1_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] PF1_MSI_CAP_NEXTPTR = 8'h00;
  parameter [11:0] PF1_PB_CAP_NEXTPTR = 12'h000;
  parameter PF1_PB_CAP_SYSTEM_ALLOCATED = "FALSE";
  parameter [3:0] PF1_PB_CAP_VER = 4'h1;
  parameter [7:0] PF1_PM_CAP_ID = 8'h01;
  parameter [7:0] PF1_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] PF1_PM_CAP_VER_ID = 3'h3;
  parameter PF1_RBAR_CAP_ENABLE = "FALSE";
  parameter [2:0] PF1_RBAR_CAP_INDEX0 = 3'h0;
  parameter [2:0] PF1_RBAR_CAP_INDEX1 = 3'h0;
  parameter [2:0] PF1_RBAR_CAP_INDEX2 = 3'h0;
  parameter [11:0] PF1_RBAR_CAP_NEXTPTR = 12'h000;
  parameter [19:0] PF1_RBAR_CAP_SIZE0 = 20'h00000;
  parameter [19:0] PF1_RBAR_CAP_SIZE1 = 20'h00000;
  parameter [19:0] PF1_RBAR_CAP_SIZE2 = 20'h00000;
  parameter [3:0] PF1_RBAR_CAP_VER = 4'h1;
  parameter [2:0] PF1_RBAR_NUM = 3'h1;
  parameter [7:0] PF1_REVISION_ID = 8'h00;
  parameter [4:0] PF1_SRIOV_BAR0_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_SRIOV_BAR0_CONTROL = 3'h4;
  parameter [4:0] PF1_SRIOV_BAR1_APERTURE_SIZE = 5'h00;
  parameter [2:0] PF1_SRIOV_BAR1_CONTROL = 3'h0;
  parameter [4:0] PF1_SRIOV_BAR2_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_SRIOV_BAR2_CONTROL = 3'h4;
  parameter [4:0] PF1_SRIOV_BAR3_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_SRIOV_BAR3_CONTROL = 3'h0;
  parameter [4:0] PF1_SRIOV_BAR4_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_SRIOV_BAR4_CONTROL = 3'h4;
  parameter [4:0] PF1_SRIOV_BAR5_APERTURE_SIZE = 5'h03;
  parameter [2:0] PF1_SRIOV_BAR5_CONTROL = 3'h0;
  parameter [15:0] PF1_SRIOV_CAP_INITIAL_VF = 16'h0000;
  parameter [11:0] PF1_SRIOV_CAP_NEXTPTR = 12'h000;
  parameter [15:0] PF1_SRIOV_CAP_TOTAL_VF = 16'h0000;
  parameter [3:0] PF1_SRIOV_CAP_VER = 4'h1;
  parameter [15:0] PF1_SRIOV_FIRST_VF_OFFSET = 16'h0000;
  parameter [15:0] PF1_SRIOV_FUNC_DEP_LINK = 16'h0000;
  parameter [31:0] PF1_SRIOV_SUPPORTED_PAGE_SIZE = 32'h00000000;
  parameter [15:0] PF1_SRIOV_VF_DEVICE_ID = 16'h0000;
  parameter [15:0] PF1_SUBSYSTEM_ID = 16'h0000;
  parameter PF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter PF1_TPHR_CAP_ENABLE = "FALSE";
  parameter PF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] PF1_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] PF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] PF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] PF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] PF1_TPHR_CAP_VER = 4'h1;
  parameter PL_DISABLE_EI_INFER_IN_L0 = "FALSE";
  parameter PL_DISABLE_GEN3_DC_BALANCE = "FALSE";
  parameter PL_DISABLE_SCRAMBLING = "FALSE";
  parameter PL_DISABLE_UPCONFIG_CAPABLE = "FALSE";
  parameter PL_EQ_ADAPT_DISABLE_COEFF_CHECK = "FALSE";
  parameter PL_EQ_ADAPT_DISABLE_PRESET_CHECK = "FALSE";
  parameter [4:0] PL_EQ_ADAPT_ITER_COUNT = 5'h02;
  parameter [1:0] PL_EQ_ADAPT_REJECT_RETRY_COUNT = 2'h1;
  parameter PL_EQ_BYPASS_PHASE23 = "FALSE";
  parameter PL_EQ_SHORT_ADAPT_PHASE = "FALSE";
  parameter [15:0] PL_LANE0_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE1_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE2_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE3_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE4_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE5_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE6_EQ_CONTROL = 16'h3F00;
  parameter [15:0] PL_LANE7_EQ_CONTROL = 16'h3F00;
  parameter [2:0] PL_LINK_CAP_MAX_LINK_SPEED = 3'h4;
  parameter [3:0] PL_LINK_CAP_MAX_LINK_WIDTH = 4'h8;
  parameter integer PL_N_FTS_COMCLK_GEN1 = 255;
  parameter integer PL_N_FTS_COMCLK_GEN2 = 255;
  parameter integer PL_N_FTS_COMCLK_GEN3 = 255;
  parameter integer PL_N_FTS_GEN1 = 255;
  parameter integer PL_N_FTS_GEN2 = 255;
  parameter integer PL_N_FTS_GEN3 = 255;
  parameter PL_SIM_FAST_LINK_TRAINING = "FALSE";
  parameter PL_UPSTREAM_FACING = "TRUE";
  parameter [15:0] PM_ASPML0S_TIMEOUT = 16'h05DC;
  parameter [19:0] PM_ASPML1_ENTRY_DELAY = 20'h00000;
  parameter PM_ENABLE_SLOT_POWER_CAPTURE = "TRUE";
  parameter [31:0] PM_L1_REENTRY_DELAY = 32'h00000000;
  parameter [19:0] PM_PME_SERVICE_TIMEOUT_DELAY = 20'h186A0;
  parameter [15:0] PM_PME_TURNOFF_ACK_DELAY = 16'h0064;
  parameter SIM_VERSION = "1.0";
  parameter integer SPARE_BIT0 = 0;
  parameter integer SPARE_BIT1 = 0;
  parameter integer SPARE_BIT2 = 0;
  parameter integer SPARE_BIT3 = 0;
  parameter integer SPARE_BIT4 = 0;
  parameter integer SPARE_BIT5 = 0;
  parameter integer SPARE_BIT6 = 0;
  parameter integer SPARE_BIT7 = 0;
  parameter integer SPARE_BIT8 = 0;
  parameter [7:0] SPARE_BYTE0 = 8'h00;
  parameter [7:0] SPARE_BYTE1 = 8'h00;
  parameter [7:0] SPARE_BYTE2 = 8'h00;
  parameter [7:0] SPARE_BYTE3 = 8'h00;
  parameter [31:0] SPARE_WORD0 = 32'h00000000;
  parameter [31:0] SPARE_WORD1 = 32'h00000000;
  parameter [31:0] SPARE_WORD2 = 32'h00000000;
  parameter [31:0] SPARE_WORD3 = 32'h00000000;
  parameter SRIOV_CAP_ENABLE = "FALSE";
  parameter [23:0] TL_COMPL_TIMEOUT_REG0 = 24'hBEBC20;
  parameter [27:0] TL_COMPL_TIMEOUT_REG1 = 28'h0000000;
  parameter [11:0] TL_CREDITS_CD = 12'h3E0;
  parameter [7:0] TL_CREDITS_CH = 8'h20;
  parameter [11:0] TL_CREDITS_NPD = 12'h028;
  parameter [7:0] TL_CREDITS_NPH = 8'h20;
  parameter [11:0] TL_CREDITS_PD = 12'h198;
  parameter [7:0] TL_CREDITS_PH = 8'h20;
  parameter TL_ENABLE_MESSAGE_RID_CHECK_ENABLE = "TRUE";
  parameter TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
  parameter TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE = "FALSE";
  parameter TL_LEGACY_MODE_ENABLE = "FALSE";
  parameter TL_PF_ENABLE_REG = "FALSE";
  parameter TL_TAG_MGMT_ENABLE = "TRUE";
  parameter [11:0] VF0_ARI_CAP_NEXTPTR = 12'h000;
  parameter [7:0] VF0_CAPABILITY_POINTER = 8'h50;
  parameter integer VF0_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF0_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF0_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF0_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF0_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF0_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF0_PM_CAP_ID = 8'h01;
  parameter [7:0] VF0_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF0_PM_CAP_VER_ID = 3'h3;
  parameter VF0_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF0_TPHR_CAP_ENABLE = "FALSE";
  parameter VF0_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF0_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF0_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF0_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF0_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF0_TPHR_CAP_VER = 4'h1;
  parameter [11:0] VF1_ARI_CAP_NEXTPTR = 12'h000;
  parameter integer VF1_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF1_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF1_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF1_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF1_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF1_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF1_PM_CAP_ID = 8'h01;
  parameter [7:0] VF1_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF1_PM_CAP_VER_ID = 3'h3;
  parameter VF1_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF1_TPHR_CAP_ENABLE = "FALSE";
  parameter VF1_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF1_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF1_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF1_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF1_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF1_TPHR_CAP_VER = 4'h1;
  parameter [11:0] VF2_ARI_CAP_NEXTPTR = 12'h000;
  parameter integer VF2_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF2_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF2_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF2_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF2_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF2_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF2_PM_CAP_ID = 8'h01;
  parameter [7:0] VF2_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF2_PM_CAP_VER_ID = 3'h3;
  parameter VF2_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF2_TPHR_CAP_ENABLE = "FALSE";
  parameter VF2_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF2_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF2_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF2_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF2_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF2_TPHR_CAP_VER = 4'h1;
  parameter [11:0] VF3_ARI_CAP_NEXTPTR = 12'h000;
  parameter integer VF3_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF3_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF3_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF3_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF3_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF3_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF3_PM_CAP_ID = 8'h01;
  parameter [7:0] VF3_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF3_PM_CAP_VER_ID = 3'h3;
  parameter VF3_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF3_TPHR_CAP_ENABLE = "FALSE";
  parameter VF3_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF3_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF3_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF3_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF3_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF3_TPHR_CAP_VER = 4'h1;
  parameter [11:0] VF4_ARI_CAP_NEXTPTR = 12'h000;
  parameter integer VF4_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF4_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF4_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF4_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF4_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF4_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF4_PM_CAP_ID = 8'h01;
  parameter [7:0] VF4_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF4_PM_CAP_VER_ID = 3'h3;
  parameter VF4_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF4_TPHR_CAP_ENABLE = "FALSE";
  parameter VF4_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF4_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF4_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF4_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF4_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF4_TPHR_CAP_VER = 4'h1;
  parameter [11:0] VF5_ARI_CAP_NEXTPTR = 12'h000;
  parameter integer VF5_MSIX_CAP_PBA_BIR = 0;
  parameter [28:0] VF5_MSIX_CAP_PBA_OFFSET = 29'h00000050;
  parameter integer VF5_MSIX_CAP_TABLE_BIR = 0;
  parameter [28:0] VF5_MSIX_CAP_TABLE_OFFSET = 29'h00000040;
  parameter [10:0] VF5_MSIX_CAP_TABLE_SIZE = 11'h000;
  parameter integer VF5_MSI_CAP_MULTIMSGCAP = 0;
  parameter [7:0] VF5_PM_CAP_ID = 8'h01;
  parameter [7:0] VF5_PM_CAP_NEXTPTR = 8'h00;
  parameter [2:0] VF5_PM_CAP_VER_ID = 3'h3;
  parameter VF5_TPHR_CAP_DEV_SPECIFIC_MODE = "TRUE";
  parameter VF5_TPHR_CAP_ENABLE = "FALSE";
  parameter VF5_TPHR_CAP_INT_VEC_MODE = "TRUE";
  parameter [11:0] VF5_TPHR_CAP_NEXTPTR = 12'h000;
  parameter [2:0] VF5_TPHR_CAP_ST_MODE_SEL = 3'h0;
  parameter [1:0] VF5_TPHR_CAP_ST_TABLE_LOC = 2'h0;
  parameter [10:0] VF5_TPHR_CAP_ST_TABLE_SIZE = 11'h000;
  parameter [3:0] VF5_TPHR_CAP_VER = 4'h1;
  
  localparam in_delay = 0;
  localparam out_delay = 0;
  localparam INCLK_DELAY = 0;
  localparam OUTCLK_DELAY = 0;

  output CFGERRCOROUT;
  output CFGERRFATALOUT;
  output CFGERRNONFATALOUT;
  output CFGEXTREADRECEIVED;
  output CFGEXTWRITERECEIVED;
  output CFGHOTRESETOUT;
  output CFGINPUTUPDATEDONE;
  output CFGINTERRUPTAOUTPUT;
  output CFGINTERRUPTBOUTPUT;
  output CFGINTERRUPTCOUTPUT;
  output CFGINTERRUPTDOUTPUT;
  output CFGINTERRUPTMSIFAIL;
  output CFGINTERRUPTMSIMASKUPDATE;
  output CFGINTERRUPTMSISENT;
  output CFGINTERRUPTMSIXFAIL;
  output CFGINTERRUPTMSIXSENT;
  output CFGINTERRUPTSENT;
  output CFGLOCALERROR;
  output CFGLTRENABLE;
  output CFGMCUPDATEDONE;
  output CFGMGMTREADWRITEDONE;
  output CFGMSGRECEIVED;
  output CFGMSGTRANSMITDONE;
  output CFGPERFUNCTIONUPDATEDONE;
  output CFGPHYLINKDOWN;
  output CFGPLSTATUSCHANGE;
  output CFGPOWERSTATECHANGEINTERRUPT;
  output CFGTPHSTTREADENABLE;
  output CFGTPHSTTWRITEENABLE;
  output DRPRDY;
  output MAXISCQTLAST;
  output MAXISCQTVALID;
  output MAXISRCTLAST;
  output MAXISRCTVALID;
  output PCIERQSEQNUMVLD;
  output PCIERQTAGVLD;
  output PIPERX0POLARITY;
  output PIPERX1POLARITY;
  output PIPERX2POLARITY;
  output PIPERX3POLARITY;
  output PIPERX4POLARITY;
  output PIPERX5POLARITY;
  output PIPERX6POLARITY;
  output PIPERX7POLARITY;
  output PIPETX0COMPLIANCE;
  output PIPETX0DATAVALID;
  output PIPETX0ELECIDLE;
  output PIPETX0STARTBLOCK;
  output PIPETX1COMPLIANCE;
  output PIPETX1DATAVALID;
  output PIPETX1ELECIDLE;
  output PIPETX1STARTBLOCK;
  output PIPETX2COMPLIANCE;
  output PIPETX2DATAVALID;
  output PIPETX2ELECIDLE;
  output PIPETX2STARTBLOCK;
  output PIPETX3COMPLIANCE;
  output PIPETX3DATAVALID;
  output PIPETX3ELECIDLE;
  output PIPETX3STARTBLOCK;
  output PIPETX4COMPLIANCE;
  output PIPETX4DATAVALID;
  output PIPETX4ELECIDLE;
  output PIPETX4STARTBLOCK;
  output PIPETX5COMPLIANCE;
  output PIPETX5DATAVALID;
  output PIPETX5ELECIDLE;
  output PIPETX5STARTBLOCK;
  output PIPETX6COMPLIANCE;
  output PIPETX6DATAVALID;
  output PIPETX6ELECIDLE;
  output PIPETX6STARTBLOCK;
  output PIPETX7COMPLIANCE;
  output PIPETX7DATAVALID;
  output PIPETX7ELECIDLE;
  output PIPETX7STARTBLOCK;
  output PIPETXDEEMPH;
  output PIPETXRCVRDET;
  output PIPETXRESET;
  output PIPETXSWING;
  output PLEQINPROGRESS;
  output [11:0] CFGFCCPLD;
  output [11:0] CFGFCNPD;
  output [11:0] CFGFCPD;
  output [11:0] CFGVFSTATUS;
  output [143:0] MIREPLAYRAMWRITEDATA;
  output [143:0] MIREQUESTRAMWRITEDATA;
  output [15:0] CFGPERFUNCSTATUSDATA;
  output [15:0] DBGDATAOUT;
  output [15:0] DRPDO;
  output [17:0] CFGVFPOWERSTATE;
  output [17:0] CFGVFTPHSTMODE;
  output [1:0] CFGDPASUBSTATECHANGE;
  output [1:0] CFGFLRINPROCESS;
  output [1:0] CFGINTERRUPTMSIENABLE;
  output [1:0] CFGINTERRUPTMSIXENABLE;
  output [1:0] CFGINTERRUPTMSIXMASK;
  output [1:0] CFGLINKPOWERSTATE;
  output [1:0] CFGOBFFENABLE;
  output [1:0] CFGPHYLINKSTATUS;
  output [1:0] CFGRCBSTATUS;
  output [1:0] CFGTPHREQUESTERENABLE;
  output [1:0] MIREPLAYRAMREADENABLE;
  output [1:0] MIREPLAYRAMWRITEENABLE;
  output [1:0] PCIERQTAGAV;
  output [1:0] PCIETFCNPDAV;
  output [1:0] PCIETFCNPHAV;
  output [1:0] PIPERX0EQCONTROL;
  output [1:0] PIPERX1EQCONTROL;
  output [1:0] PIPERX2EQCONTROL;
  output [1:0] PIPERX3EQCONTROL;
  output [1:0] PIPERX4EQCONTROL;
  output [1:0] PIPERX5EQCONTROL;
  output [1:0] PIPERX6EQCONTROL;
  output [1:0] PIPERX7EQCONTROL;
  output [1:0] PIPETX0CHARISK;
  output [1:0] PIPETX0EQCONTROL;
  output [1:0] PIPETX0POWERDOWN;
  output [1:0] PIPETX0SYNCHEADER;
  output [1:0] PIPETX1CHARISK;
  output [1:0] PIPETX1EQCONTROL;
  output [1:0] PIPETX1POWERDOWN;
  output [1:0] PIPETX1SYNCHEADER;
  output [1:0] PIPETX2CHARISK;
  output [1:0] PIPETX2EQCONTROL;
  output [1:0] PIPETX2POWERDOWN;
  output [1:0] PIPETX2SYNCHEADER;
  output [1:0] PIPETX3CHARISK;
  output [1:0] PIPETX3EQCONTROL;
  output [1:0] PIPETX3POWERDOWN;
  output [1:0] PIPETX3SYNCHEADER;
  output [1:0] PIPETX4CHARISK;
  output [1:0] PIPETX4EQCONTROL;
  output [1:0] PIPETX4POWERDOWN;
  output [1:0] PIPETX4SYNCHEADER;
  output [1:0] PIPETX5CHARISK;
  output [1:0] PIPETX5EQCONTROL;
  output [1:0] PIPETX5POWERDOWN;
  output [1:0] PIPETX5SYNCHEADER;
  output [1:0] PIPETX6CHARISK;
  output [1:0] PIPETX6EQCONTROL;
  output [1:0] PIPETX6POWERDOWN;
  output [1:0] PIPETX6SYNCHEADER;
  output [1:0] PIPETX7CHARISK;
  output [1:0] PIPETX7EQCONTROL;
  output [1:0] PIPETX7POWERDOWN;
  output [1:0] PIPETX7SYNCHEADER;
  output [1:0] PIPETXRATE;
  output [1:0] PLEQPHASE;
  output [255:0] MAXISCQTDATA;
  output [255:0] MAXISRCTDATA;
  output [2:0] CFGCURRENTSPEED;
  output [2:0] CFGMAXPAYLOAD;
  output [2:0] CFGMAXREADREQ;
  output [2:0] CFGTPHFUNCTIONNUM;
  output [2:0] PIPERX0EQPRESET;
  output [2:0] PIPERX1EQPRESET;
  output [2:0] PIPERX2EQPRESET;
  output [2:0] PIPERX3EQPRESET;
  output [2:0] PIPERX4EQPRESET;
  output [2:0] PIPERX5EQPRESET;
  output [2:0] PIPERX6EQPRESET;
  output [2:0] PIPERX7EQPRESET;
  output [2:0] PIPETXMARGIN;
  output [31:0] CFGEXTWRITEDATA;
  output [31:0] CFGINTERRUPTMSIDATA;
  output [31:0] CFGMGMTREADDATA;
  output [31:0] CFGTPHSTTWRITEDATA;
  output [31:0] PIPETX0DATA;
  output [31:0] PIPETX1DATA;
  output [31:0] PIPETX2DATA;
  output [31:0] PIPETX3DATA;
  output [31:0] PIPETX4DATA;
  output [31:0] PIPETX5DATA;
  output [31:0] PIPETX6DATA;
  output [31:0] PIPETX7DATA;
  output [3:0] CFGEXTWRITEBYTEENABLE;
  output [3:0] CFGNEGOTIATEDWIDTH;
  output [3:0] CFGTPHSTTWRITEBYTEVALID;
  output [3:0] MICOMPLETIONRAMREADENABLEL;
  output [3:0] MICOMPLETIONRAMREADENABLEU;
  output [3:0] MICOMPLETIONRAMWRITEENABLEL;
  output [3:0] MICOMPLETIONRAMWRITEENABLEU;
  output [3:0] MIREQUESTRAMREADENABLE;
  output [3:0] MIREQUESTRAMWRITEENABLE;
  output [3:0] PCIERQSEQNUM;
  output [3:0] PIPERX0EQLPTXPRESET;
  output [3:0] PIPERX1EQLPTXPRESET;
  output [3:0] PIPERX2EQLPTXPRESET;
  output [3:0] PIPERX3EQLPTXPRESET;
  output [3:0] PIPERX4EQLPTXPRESET;
  output [3:0] PIPERX5EQLPTXPRESET;
  output [3:0] PIPERX6EQLPTXPRESET;
  output [3:0] PIPERX7EQLPTXPRESET;
  output [3:0] PIPETX0EQPRESET;
  output [3:0] PIPETX1EQPRESET;
  output [3:0] PIPETX2EQPRESET;
  output [3:0] PIPETX3EQPRESET;
  output [3:0] PIPETX4EQPRESET;
  output [3:0] PIPETX5EQPRESET;
  output [3:0] PIPETX6EQPRESET;
  output [3:0] PIPETX7EQPRESET;
  output [3:0] SAXISCCTREADY;
  output [3:0] SAXISRQTREADY;
  output [4:0] CFGMSGRECEIVEDTYPE;
  output [4:0] CFGTPHSTTADDRESS;
  output [5:0] CFGFUNCTIONPOWERSTATE;
  output [5:0] CFGINTERRUPTMSIMMENABLE;
  output [5:0] CFGINTERRUPTMSIVFENABLE;
  output [5:0] CFGINTERRUPTMSIXVFENABLE;
  output [5:0] CFGINTERRUPTMSIXVFMASK;
  output [5:0] CFGLTSSMSTATE;
  output [5:0] CFGTPHSTMODE;
  output [5:0] CFGVFFLRINPROCESS;
  output [5:0] CFGVFTPHREQUESTERENABLE;
  output [5:0] PCIECQNPREQCOUNT;
  output [5:0] PCIERQTAG;
  output [5:0] PIPERX0EQLPLFFS;
  output [5:0] PIPERX1EQLPLFFS;
  output [5:0] PIPERX2EQLPLFFS;
  output [5:0] PIPERX3EQLPLFFS;
  output [5:0] PIPERX4EQLPLFFS;
  output [5:0] PIPERX5EQLPLFFS;
  output [5:0] PIPERX6EQLPLFFS;
  output [5:0] PIPERX7EQLPLFFS;
  output [5:0] PIPETX0EQDEEMPH;
  output [5:0] PIPETX1EQDEEMPH;
  output [5:0] PIPETX2EQDEEMPH;
  output [5:0] PIPETX3EQDEEMPH;
  output [5:0] PIPETX4EQDEEMPH;
  output [5:0] PIPETX5EQDEEMPH;
  output [5:0] PIPETX6EQDEEMPH;
  output [5:0] PIPETX7EQDEEMPH;
  output [71:0] MICOMPLETIONRAMWRITEDATAL;
  output [71:0] MICOMPLETIONRAMWRITEDATAU;
  output [74:0] MAXISRCTUSER;
  output [7:0] CFGEXTFUNCTIONNUMBER;
  output [7:0] CFGFCCPLH;
  output [7:0] CFGFCNPH;
  output [7:0] CFGFCPH;
  output [7:0] CFGFUNCTIONSTATUS;
  output [7:0] CFGMSGRECEIVEDDATA;
  output [7:0] MAXISCQTKEEP;
  output [7:0] MAXISRCTKEEP;
  output [7:0] PLGEN3PCSRXSLIDE;
  output [84:0] MAXISCQTUSER;
  output [8:0] MIREPLAYRAMADDRESS;
  output [8:0] MIREQUESTRAMREADADDRESSA;
  output [8:0] MIREQUESTRAMREADADDRESSB;
  output [8:0] MIREQUESTRAMWRITEADDRESSA;
  output [8:0] MIREQUESTRAMWRITEADDRESSB;
  output [9:0] CFGEXTREGISTERNUMBER;
  output [9:0] MICOMPLETIONRAMREADADDRESSAL;
  output [9:0] MICOMPLETIONRAMREADADDRESSAU;
  output [9:0] MICOMPLETIONRAMREADADDRESSBL;
  output [9:0] MICOMPLETIONRAMREADADDRESSBU;
  output [9:0] MICOMPLETIONRAMWRITEADDRESSAL;
  output [9:0] MICOMPLETIONRAMWRITEADDRESSAU;
  output [9:0] MICOMPLETIONRAMWRITEADDRESSBL;
  output [9:0] MICOMPLETIONRAMWRITEADDRESSBU;

  input CFGCONFIGSPACEENABLE;
  input CFGERRCORIN;
  input CFGERRUNCORIN;
  input CFGEXTREADDATAVALID;
  input CFGHOTRESETIN;
  input CFGINPUTUPDATEREQUEST;
  input CFGINTERRUPTMSITPHPRESENT;
  input CFGINTERRUPTMSIXINT;
  input CFGLINKTRAININGENABLE;
  input CFGMCUPDATEREQUEST;
  input CFGMGMTREAD;
  input CFGMGMTTYPE1CFGREGACCESS;
  input CFGMGMTWRITE;
  input CFGMSGTRANSMIT;
  input CFGPERFUNCTIONOUTPUTREQUEST;
  input CFGPOWERSTATECHANGEACK;
  input CFGREQPMTRANSITIONL23READY;
  input CFGTPHSTTREADDATAVALID;
  input CORECLK;
  input CORECLKMICOMPLETIONRAML;
  input CORECLKMICOMPLETIONRAMU;
  input CORECLKMIREPLAYRAM;
  input CORECLKMIREQUESTRAM;
  input DRPCLK;
  input DRPEN;
  input DRPWE;
  input MGMTRESETN;
  input MGMTSTICKYRESETN;
  input PCIECQNPREQ;
  input PIPECLK;
  input PIPERESETN;
  input PIPERX0DATAVALID;
  input PIPERX0ELECIDLE;
  input PIPERX0EQDONE;
  input PIPERX0EQLPADAPTDONE;
  input PIPERX0EQLPLFFSSEL;
  input PIPERX0PHYSTATUS;
  input PIPERX0STARTBLOCK;
  input PIPERX0VALID;
  input PIPERX1DATAVALID;
  input PIPERX1ELECIDLE;
  input PIPERX1EQDONE;
  input PIPERX1EQLPADAPTDONE;
  input PIPERX1EQLPLFFSSEL;
  input PIPERX1PHYSTATUS;
  input PIPERX1STARTBLOCK;
  input PIPERX1VALID;
  input PIPERX2DATAVALID;
  input PIPERX2ELECIDLE;
  input PIPERX2EQDONE;
  input PIPERX2EQLPADAPTDONE;
  input PIPERX2EQLPLFFSSEL;
  input PIPERX2PHYSTATUS;
  input PIPERX2STARTBLOCK;
  input PIPERX2VALID;
  input PIPERX3DATAVALID;
  input PIPERX3ELECIDLE;
  input PIPERX3EQDONE;
  input PIPERX3EQLPADAPTDONE;
  input PIPERX3EQLPLFFSSEL;
  input PIPERX3PHYSTATUS;
  input PIPERX3STARTBLOCK;
  input PIPERX3VALID;
  input PIPERX4DATAVALID;
  input PIPERX4ELECIDLE;
  input PIPERX4EQDONE;
  input PIPERX4EQLPADAPTDONE;
  input PIPERX4EQLPLFFSSEL;
  input PIPERX4PHYSTATUS;
  input PIPERX4STARTBLOCK;
  input PIPERX4VALID;
  input PIPERX5DATAVALID;
  input PIPERX5ELECIDLE;
  input PIPERX5EQDONE;
  input PIPERX5EQLPADAPTDONE;
  input PIPERX5EQLPLFFSSEL;
  input PIPERX5PHYSTATUS;
  input PIPERX5STARTBLOCK;
  input PIPERX5VALID;
  input PIPERX6DATAVALID;
  input PIPERX6ELECIDLE;
  input PIPERX6EQDONE;
  input PIPERX6EQLPADAPTDONE;
  input PIPERX6EQLPLFFSSEL;
  input PIPERX6PHYSTATUS;
  input PIPERX6STARTBLOCK;
  input PIPERX6VALID;
  input PIPERX7DATAVALID;
  input PIPERX7ELECIDLE;
  input PIPERX7EQDONE;
  input PIPERX7EQLPADAPTDONE;
  input PIPERX7EQLPLFFSSEL;
  input PIPERX7PHYSTATUS;
  input PIPERX7STARTBLOCK;
  input PIPERX7VALID;
  input PIPETX0EQDONE;
  input PIPETX1EQDONE;
  input PIPETX2EQDONE;
  input PIPETX3EQDONE;
  input PIPETX4EQDONE;
  input PIPETX5EQDONE;
  input PIPETX6EQDONE;
  input PIPETX7EQDONE;
  input PLDISABLESCRAMBLER;
  input PLEQRESETEIEOSCOUNT;
  input PLGEN3PCSDISABLE;
  input RECCLK;
  input RESETN;
  input SAXISCCTLAST;
  input SAXISCCTVALID;
  input SAXISRQTLAST;
  input SAXISRQTVALID;
  input USERCLK;
  input [10:0] DRPADDR;
  input [143:0] MICOMPLETIONRAMREADDATA;
  input [143:0] MIREPLAYRAMREADDATA;
  input [143:0] MIREQUESTRAMREADDATA;
  input [15:0] CFGDEVID;
  input [15:0] CFGSUBSYSID;
  input [15:0] CFGSUBSYSVENDID;
  input [15:0] CFGVENDID;
  input [15:0] DRPDI;
  input [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET;
  input [17:0] PIPETX0EQCOEFF;
  input [17:0] PIPETX1EQCOEFF;
  input [17:0] PIPETX2EQCOEFF;
  input [17:0] PIPETX3EQCOEFF;
  input [17:0] PIPETX4EQCOEFF;
  input [17:0] PIPETX5EQCOEFF;
  input [17:0] PIPETX6EQCOEFF;
  input [17:0] PIPETX7EQCOEFF;
  input [18:0] CFGMGMTADDR;
  input [1:0] CFGFLRDONE;
  input [1:0] CFGINTERRUPTMSITPHTYPE;
  input [1:0] CFGINTERRUPTPENDING;
  input [1:0] PIPERX0CHARISK;
  input [1:0] PIPERX0SYNCHEADER;
  input [1:0] PIPERX1CHARISK;
  input [1:0] PIPERX1SYNCHEADER;
  input [1:0] PIPERX2CHARISK;
  input [1:0] PIPERX2SYNCHEADER;
  input [1:0] PIPERX3CHARISK;
  input [1:0] PIPERX3SYNCHEADER;
  input [1:0] PIPERX4CHARISK;
  input [1:0] PIPERX4SYNCHEADER;
  input [1:0] PIPERX5CHARISK;
  input [1:0] PIPERX5SYNCHEADER;
  input [1:0] PIPERX6CHARISK;
  input [1:0] PIPERX6SYNCHEADER;
  input [1:0] PIPERX7CHARISK;
  input [1:0] PIPERX7SYNCHEADER;
  input [21:0] MAXISCQTREADY;
  input [21:0] MAXISRCTREADY;
  input [255:0] SAXISCCTDATA;
  input [255:0] SAXISRQTDATA;
  input [2:0] CFGDSFUNCTIONNUMBER;
  input [2:0] CFGFCSEL;
  input [2:0] CFGINTERRUPTMSIATTR;
  input [2:0] CFGINTERRUPTMSIFUNCTIONNUMBER;
  input [2:0] CFGMSGTRANSMITTYPE;
  input [2:0] CFGPERFUNCSTATUSCONTROL;
  input [2:0] CFGPERFUNCTIONNUMBER;
  input [2:0] PIPERX0STATUS;
  input [2:0] PIPERX1STATUS;
  input [2:0] PIPERX2STATUS;
  input [2:0] PIPERX3STATUS;
  input [2:0] PIPERX4STATUS;
  input [2:0] PIPERX5STATUS;
  input [2:0] PIPERX6STATUS;
  input [2:0] PIPERX7STATUS;
  input [31:0] CFGEXTREADDATA;
  input [31:0] CFGINTERRUPTMSIINT;
  input [31:0] CFGINTERRUPTMSIXDATA;
  input [31:0] CFGMGMTWRITEDATA;
  input [31:0] CFGMSGTRANSMITDATA;
  input [31:0] CFGTPHSTTREADDATA;
  input [31:0] PIPERX0DATA;
  input [31:0] PIPERX1DATA;
  input [31:0] PIPERX2DATA;
  input [31:0] PIPERX3DATA;
  input [31:0] PIPERX4DATA;
  input [31:0] PIPERX5DATA;
  input [31:0] PIPERX6DATA;
  input [31:0] PIPERX7DATA;
  input [32:0] SAXISCCTUSER;
  input [3:0] CFGINTERRUPTINT;
  input [3:0] CFGINTERRUPTMSISELECT;
  input [3:0] CFGMGMTBYTEENABLE;
  input [4:0] CFGDSDEVICENUMBER;
  input [59:0] SAXISRQTUSER;
  input [5:0] CFGVFFLRDONE;
  input [5:0] PIPEEQFS;
  input [5:0] PIPEEQLF;
  input [63:0] CFGDSN;
  input [63:0] CFGINTERRUPTMSIPENDINGSTATUS;
  input [63:0] CFGINTERRUPTMSIXADDRESS;
  input [7:0] CFGDSBUSNUMBER;
  input [7:0] CFGDSPORTNUMBER;
  input [7:0] CFGREVID;
  input [7:0] PLGEN3PCSRXSYNCDONE;
  input [7:0] SAXISCCTKEEP;
  input [7:0] SAXISRQTKEEP;
  input [8:0] CFGINTERRUPTMSITPHSTTAG;

  reg SIM_VERSION_BINARY;
  reg [0:0] ARI_CAP_ENABLE_BINARY;
  reg [0:0] AXISTEN_IF_CC_ALIGNMENT_MODE_BINARY;
  reg [0:0] AXISTEN_IF_CC_PARITY_CHK_BINARY;
  reg [0:0] AXISTEN_IF_CQ_ALIGNMENT_MODE_BINARY;
  reg [0:0] AXISTEN_IF_ENABLE_CLIENT_TAG_BINARY;
  reg [0:0] AXISTEN_IF_ENABLE_RX_MSG_INTFC_BINARY;
  reg [0:0] AXISTEN_IF_RC_ALIGNMENT_MODE_BINARY;
  reg [0:0] AXISTEN_IF_RC_STRADDLE_BINARY;
  reg [0:0] AXISTEN_IF_RQ_ALIGNMENT_MODE_BINARY;
  reg [0:0] AXISTEN_IF_RQ_PARITY_CHK_BINARY;
  reg [0:0] CRM_CORE_CLK_FREQ_500_BINARY;
  reg [0:0] GEN3_PCS_RX_ELECIDLE_INTERNAL_BINARY;
  reg [0:0] LL_ACK_TIMEOUT_EN_BINARY;
  reg [0:0] LL_CPL_FC_UPDATE_TIMER_OVERRIDE_BINARY;
  reg [0:0] LL_FC_UPDATE_TIMER_OVERRIDE_BINARY;
  reg [0:0] LL_NP_FC_UPDATE_TIMER_OVERRIDE_BINARY;
  reg [0:0] LL_P_FC_UPDATE_TIMER_OVERRIDE_BINARY;
  reg [0:0] LL_REPLAY_TIMEOUT_EN_BINARY;
  reg [0:0] LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_BINARY;
  reg [0:0] LTR_TX_MESSAGE_ON_LTR_ENABLE_BINARY;
  reg [0:0] PF0_AER_CAP_ECRC_CHECK_CAPABLE_BINARY;
  reg [0:0] PF0_AER_CAP_ECRC_GEN_CAPABLE_BINARY;
  reg [0:0] PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_BINARY;
  reg [0:0] PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_BINARY;
  reg [0:0] PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_BINARY;
  reg [0:0] PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_BINARY;
  reg [0:0] PF0_DEV_CAP2_LTR_SUPPORT_BINARY;
  reg [0:0] PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_BINARY;
  reg [0:0] PF0_DEV_CAP_EXT_TAG_SUPPORTED_BINARY;
  reg [0:0] PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_BINARY;
  reg [0:0] PF0_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY;
  reg [0:0] PF0_EXPANSION_ROM_ENABLE_BINARY;
  reg [0:0] PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_BINARY;
  reg [0:0] PF0_PB_CAP_SYSTEM_ALLOCATED_BINARY;
  reg [0:0] PF0_PM_CAP_PMESUPPORT_D0_BINARY;
  reg [0:0] PF0_PM_CAP_PMESUPPORT_D1_BINARY;
  reg [0:0] PF0_PM_CAP_PMESUPPORT_D3HOT_BINARY;
  reg [0:0] PF0_PM_CAP_SUPP_D1_STATE_BINARY;
  reg [0:0] PF0_PM_CSR_NOSOFTRESET_BINARY;
  reg [0:0] PF0_RBAR_CAP_ENABLE_BINARY;
  reg [0:0] PF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] PF0_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] PF0_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] PF1_AER_CAP_ECRC_CHECK_CAPABLE_BINARY;
  reg [0:0] PF1_AER_CAP_ECRC_GEN_CAPABLE_BINARY;
  reg [0:0] PF1_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY;
  reg [0:0] PF1_EXPANSION_ROM_ENABLE_BINARY;
  reg [0:0] PF1_PB_CAP_SYSTEM_ALLOCATED_BINARY;
  reg [0:0] PF1_RBAR_CAP_ENABLE_BINARY;
  reg [0:0] PF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] PF1_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] PF1_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] PL_DISABLE_EI_INFER_IN_L0_BINARY;
  reg [0:0] PL_DISABLE_GEN3_DC_BALANCE_BINARY;
  reg [0:0] PL_DISABLE_SCRAMBLING_BINARY;
  reg [0:0] PL_DISABLE_UPCONFIG_CAPABLE_BINARY;
  reg [0:0] PL_EQ_ADAPT_DISABLE_COEFF_CHECK_BINARY;
  reg [0:0] PL_EQ_ADAPT_DISABLE_PRESET_CHECK_BINARY;
  reg [0:0] PL_EQ_BYPASS_PHASE23_BINARY;
  reg [0:0] PL_EQ_SHORT_ADAPT_PHASE_BINARY;
  reg [0:0] PL_SIM_FAST_LINK_TRAINING_BINARY;
  reg [0:0] PL_UPSTREAM_FACING_BINARY;
  reg [0:0] PM_ENABLE_SLOT_POWER_CAPTURE_BINARY;
  reg [0:0] SPARE_BIT0_BINARY;
  reg [0:0] SPARE_BIT1_BINARY;
  reg [0:0] SPARE_BIT2_BINARY;
  reg [0:0] SPARE_BIT3_BINARY;
  reg [0:0] SPARE_BIT4_BINARY;
  reg [0:0] SPARE_BIT5_BINARY;
  reg [0:0] SPARE_BIT6_BINARY;
  reg [0:0] SPARE_BIT7_BINARY;
  reg [0:0] SPARE_BIT8_BINARY;
  reg [0:0] SRIOV_CAP_ENABLE_BINARY;
  reg [0:0] TL_ENABLE_MESSAGE_RID_CHECK_ENABLE_BINARY;
  reg [0:0] TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_BINARY;
  reg [0:0] TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE_BINARY;
  reg [0:0] TL_LEGACY_MODE_ENABLE_BINARY;
  reg [0:0] TL_PF_ENABLE_REG_BINARY;
  reg [0:0] TL_TAG_MGMT_ENABLE_BINARY;
  reg [0:0] VF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF0_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF0_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] VF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF1_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF1_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] VF2_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF2_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF2_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] VF3_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF3_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF3_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] VF4_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF4_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF4_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [0:0] VF5_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY;
  reg [0:0] VF5_TPHR_CAP_ENABLE_BINARY;
  reg [0:0] VF5_TPHR_CAP_INT_VEC_MODE_BINARY;
  reg [1:0] LL_ACK_TIMEOUT_FUNC_BINARY;
  reg [1:0] LL_REPLAY_TIMEOUT_FUNC_BINARY;
  reg [1:0] PF0_LINK_CAP_ASPM_SUPPORT_BINARY;
  reg [2:0] PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_BINARY;
  reg [2:0] PF0_DEV_CAP_ENDPOINT_L1_LATENCY_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_BINARY;
  reg [2:0] PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_BINARY;
  reg [2:0] PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_BINARY;
  reg [2:0] PF0_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] PF0_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] PF0_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] PF1_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] PF1_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] PF1_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF0_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF0_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF0_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF1_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF1_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF1_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF2_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF2_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF2_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF3_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF3_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF3_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF4_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF4_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF4_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [2:0] VF5_MSIX_CAP_PBA_BIR_BINARY;
  reg [2:0] VF5_MSIX_CAP_TABLE_BIR_BINARY;
  reg [2:0] VF5_MSI_CAP_MULTIMSGCAP_BINARY;
  reg [7:0] PL_N_FTS_COMCLK_GEN1_BINARY;
  reg [7:0] PL_N_FTS_COMCLK_GEN2_BINARY;
  reg [7:0] PL_N_FTS_COMCLK_GEN3_BINARY;
  reg [7:0] PL_N_FTS_GEN1_BINARY;
  reg [7:0] PL_N_FTS_GEN2_BINARY;
  reg [7:0] PL_N_FTS_GEN3_BINARY;

  reg notifier;

  wire CFGERRCOROUT_OUT;
  wire CFGERRFATALOUT_OUT;
  wire CFGERRNONFATALOUT_OUT;
  wire CFGEXTREADRECEIVED_OUT;
  wire CFGEXTWRITERECEIVED_OUT;
  wire CFGHOTRESETOUT_OUT;
  wire CFGINPUTUPDATEDONE_OUT;
  wire CFGINTERRUPTAOUTPUT_OUT;
  wire CFGINTERRUPTBOUTPUT_OUT;
  wire CFGINTERRUPTCOUTPUT_OUT;
  wire CFGINTERRUPTDOUTPUT_OUT;
  wire CFGINTERRUPTMSIFAIL_OUT;
  wire CFGINTERRUPTMSIMASKUPDATE_OUT;
  wire CFGINTERRUPTMSISENT_OUT;
  wire CFGINTERRUPTMSIXFAIL_OUT;
  wire CFGINTERRUPTMSIXSENT_OUT;
  wire CFGINTERRUPTSENT_OUT;
  wire CFGLOCALERROR_OUT;
  wire CFGLTRENABLE_OUT;
  wire CFGMCUPDATEDONE_OUT;
  wire CFGMGMTREADWRITEDONE_OUT;
  wire CFGMSGRECEIVED_OUT;
  wire CFGMSGTRANSMITDONE_OUT;
  wire CFGPERFUNCTIONUPDATEDONE_OUT;
  wire CFGPHYLINKDOWN_OUT;
  wire CFGPLSTATUSCHANGE_OUT;
  wire CFGPOWERSTATECHANGEINTERRUPT_OUT;
  wire CFGTPHSTTREADENABLE_OUT;
  wire CFGTPHSTTWRITEENABLE_OUT;
  wire DRPRDY_OUT;
  wire MAXISCQTLAST_OUT;
  wire MAXISCQTVALID_OUT;
  wire MAXISRCTLAST_OUT;
  wire MAXISRCTVALID_OUT;
  wire PCIERQSEQNUMVLD_OUT;
  wire PCIERQTAGVLD_OUT;
  wire PIPERX0POLARITY_OUT;
  wire PIPERX1POLARITY_OUT;
  wire PIPERX2POLARITY_OUT;
  wire PIPERX3POLARITY_OUT;
  wire PIPERX4POLARITY_OUT;
  wire PIPERX5POLARITY_OUT;
  wire PIPERX6POLARITY_OUT;
  wire PIPERX7POLARITY_OUT;
  wire PIPETX0COMPLIANCE_OUT;
  wire PIPETX0DATAVALID_OUT;
  wire PIPETX0ELECIDLE_OUT;
  wire PIPETX0STARTBLOCK_OUT;
  wire PIPETX1COMPLIANCE_OUT;
  wire PIPETX1DATAVALID_OUT;
  wire PIPETX1ELECIDLE_OUT;
  wire PIPETX1STARTBLOCK_OUT;
  wire PIPETX2COMPLIANCE_OUT;
  wire PIPETX2DATAVALID_OUT;
  wire PIPETX2ELECIDLE_OUT;
  wire PIPETX2STARTBLOCK_OUT;
  wire PIPETX3COMPLIANCE_OUT;
  wire PIPETX3DATAVALID_OUT;
  wire PIPETX3ELECIDLE_OUT;
  wire PIPETX3STARTBLOCK_OUT;
  wire PIPETX4COMPLIANCE_OUT;
  wire PIPETX4DATAVALID_OUT;
  wire PIPETX4ELECIDLE_OUT;
  wire PIPETX4STARTBLOCK_OUT;
  wire PIPETX5COMPLIANCE_OUT;
  wire PIPETX5DATAVALID_OUT;
  wire PIPETX5ELECIDLE_OUT;
  wire PIPETX5STARTBLOCK_OUT;
  wire PIPETX6COMPLIANCE_OUT;
  wire PIPETX6DATAVALID_OUT;
  wire PIPETX6ELECIDLE_OUT;
  wire PIPETX6STARTBLOCK_OUT;
  wire PIPETX7COMPLIANCE_OUT;
  wire PIPETX7DATAVALID_OUT;
  wire PIPETX7ELECIDLE_OUT;
  wire PIPETX7STARTBLOCK_OUT;
  wire PIPETXDEEMPH_OUT;
  wire PIPETXRCVRDET_OUT;
  wire PIPETXRESET_OUT;
  wire PIPETXSWING_OUT;
  wire PLEQINPROGRESS_OUT;
  wire [11:0] CFGFCCPLD_OUT;
  wire [11:0] CFGFCNPD_OUT;
  wire [11:0] CFGFCPD_OUT;
  wire [11:0] CFGVFSTATUS_OUT;
  wire [143:0] MIREPLAYRAMWRITEDATA_OUT;
  wire [143:0] MIREQUESTRAMWRITEDATA_OUT;
  wire [15:0] CFGPERFUNCSTATUSDATA_OUT;
  wire [15:0] DBGDATAOUT_OUT;
  wire [15:0] DRPDO_OUT;
  wire [17:0] CFGVFPOWERSTATE_OUT;
  wire [17:0] CFGVFTPHSTMODE_OUT;
  wire [1:0] CFGDPASUBSTATECHANGE_OUT;
  wire [1:0] CFGFLRINPROCESS_OUT;
  wire [1:0] CFGINTERRUPTMSIENABLE_OUT;
  wire [1:0] CFGINTERRUPTMSIXENABLE_OUT;
  wire [1:0] CFGINTERRUPTMSIXMASK_OUT;
  wire [1:0] CFGLINKPOWERSTATE_OUT;
  wire [1:0] CFGOBFFENABLE_OUT;
  wire [1:0] CFGPHYLINKSTATUS_OUT;
  wire [1:0] CFGRCBSTATUS_OUT;
  wire [1:0] CFGTPHREQUESTERENABLE_OUT;
  wire [1:0] MIREPLAYRAMREADENABLE_OUT;
  wire [1:0] MIREPLAYRAMWRITEENABLE_OUT;
  wire [1:0] PCIERQTAGAV_OUT;
  wire [1:0] PCIETFCNPDAV_OUT;
  wire [1:0] PCIETFCNPHAV_OUT;
  wire [1:0] PIPERX0EQCONTROL_OUT;
  wire [1:0] PIPERX1EQCONTROL_OUT;
  wire [1:0] PIPERX2EQCONTROL_OUT;
  wire [1:0] PIPERX3EQCONTROL_OUT;
  wire [1:0] PIPERX4EQCONTROL_OUT;
  wire [1:0] PIPERX5EQCONTROL_OUT;
  wire [1:0] PIPERX6EQCONTROL_OUT;
  wire [1:0] PIPERX7EQCONTROL_OUT;
  wire [1:0] PIPETX0CHARISK_OUT;
  wire [1:0] PIPETX0EQCONTROL_OUT;
  wire [1:0] PIPETX0POWERDOWN_OUT;
  wire [1:0] PIPETX0SYNCHEADER_OUT;
  wire [1:0] PIPETX1CHARISK_OUT;
  wire [1:0] PIPETX1EQCONTROL_OUT;
  wire [1:0] PIPETX1POWERDOWN_OUT;
  wire [1:0] PIPETX1SYNCHEADER_OUT;
  wire [1:0] PIPETX2CHARISK_OUT;
  wire [1:0] PIPETX2EQCONTROL_OUT;
  wire [1:0] PIPETX2POWERDOWN_OUT;
  wire [1:0] PIPETX2SYNCHEADER_OUT;
  wire [1:0] PIPETX3CHARISK_OUT;
  wire [1:0] PIPETX3EQCONTROL_OUT;
  wire [1:0] PIPETX3POWERDOWN_OUT;
  wire [1:0] PIPETX3SYNCHEADER_OUT;
  wire [1:0] PIPETX4CHARISK_OUT;
  wire [1:0] PIPETX4EQCONTROL_OUT;
  wire [1:0] PIPETX4POWERDOWN_OUT;
  wire [1:0] PIPETX4SYNCHEADER_OUT;
  wire [1:0] PIPETX5CHARISK_OUT;
  wire [1:0] PIPETX5EQCONTROL_OUT;
  wire [1:0] PIPETX5POWERDOWN_OUT;
  wire [1:0] PIPETX5SYNCHEADER_OUT;
  wire [1:0] PIPETX6CHARISK_OUT;
  wire [1:0] PIPETX6EQCONTROL_OUT;
  wire [1:0] PIPETX6POWERDOWN_OUT;
  wire [1:0] PIPETX6SYNCHEADER_OUT;
  wire [1:0] PIPETX7CHARISK_OUT;
  wire [1:0] PIPETX7EQCONTROL_OUT;
  wire [1:0] PIPETX7POWERDOWN_OUT;
  wire [1:0] PIPETX7SYNCHEADER_OUT;
  wire [1:0] PIPETXRATE_OUT;
  wire [1:0] PLEQPHASE_OUT;
  wire [255:0] MAXISCQTDATA_OUT;
  wire [255:0] MAXISRCTDATA_OUT;
  wire [2:0] CFGCURRENTSPEED_OUT;
  wire [2:0] CFGMAXPAYLOAD_OUT;
  wire [2:0] CFGMAXREADREQ_OUT;
  wire [2:0] CFGTPHFUNCTIONNUM_OUT;
  wire [2:0] PIPERX0EQPRESET_OUT;
  wire [2:0] PIPERX1EQPRESET_OUT;
  wire [2:0] PIPERX2EQPRESET_OUT;
  wire [2:0] PIPERX3EQPRESET_OUT;
  wire [2:0] PIPERX4EQPRESET_OUT;
  wire [2:0] PIPERX5EQPRESET_OUT;
  wire [2:0] PIPERX6EQPRESET_OUT;
  wire [2:0] PIPERX7EQPRESET_OUT;
  wire [2:0] PIPETXMARGIN_OUT;
  wire [31:0] CFGEXTWRITEDATA_OUT;
  wire [31:0] CFGINTERRUPTMSIDATA_OUT;
  wire [31:0] CFGMGMTREADDATA_OUT;
  wire [31:0] CFGTPHSTTWRITEDATA_OUT;
  wire [31:0] PIPETX0DATA_OUT;
  wire [31:0] PIPETX1DATA_OUT;
  wire [31:0] PIPETX2DATA_OUT;
  wire [31:0] PIPETX3DATA_OUT;
  wire [31:0] PIPETX4DATA_OUT;
  wire [31:0] PIPETX5DATA_OUT;
  wire [31:0] PIPETX6DATA_OUT;
  wire [31:0] PIPETX7DATA_OUT;
  wire [3:0] CFGEXTWRITEBYTEENABLE_OUT;
  wire [3:0] CFGNEGOTIATEDWIDTH_OUT;
  wire [3:0] CFGTPHSTTWRITEBYTEVALID_OUT;
  wire [3:0] MICOMPLETIONRAMREADENABLEL_OUT;
  wire [3:0] MICOMPLETIONRAMREADENABLEU_OUT;
  wire [3:0] MICOMPLETIONRAMWRITEENABLEL_OUT;
  wire [3:0] MICOMPLETIONRAMWRITEENABLEU_OUT;
  wire [3:0] MIREQUESTRAMREADENABLE_OUT;
  wire [3:0] MIREQUESTRAMWRITEENABLE_OUT;
  wire [3:0] PCIERQSEQNUM_OUT;
  wire [3:0] PIPERX0EQLPTXPRESET_OUT;
  wire [3:0] PIPERX1EQLPTXPRESET_OUT;
  wire [3:0] PIPERX2EQLPTXPRESET_OUT;
  wire [3:0] PIPERX3EQLPTXPRESET_OUT;
  wire [3:0] PIPERX4EQLPTXPRESET_OUT;
  wire [3:0] PIPERX5EQLPTXPRESET_OUT;
  wire [3:0] PIPERX6EQLPTXPRESET_OUT;
  wire [3:0] PIPERX7EQLPTXPRESET_OUT;
  wire [3:0] PIPETX0EQPRESET_OUT;
  wire [3:0] PIPETX1EQPRESET_OUT;
  wire [3:0] PIPETX2EQPRESET_OUT;
  wire [3:0] PIPETX3EQPRESET_OUT;
  wire [3:0] PIPETX4EQPRESET_OUT;
  wire [3:0] PIPETX5EQPRESET_OUT;
  wire [3:0] PIPETX6EQPRESET_OUT;
  wire [3:0] PIPETX7EQPRESET_OUT;
  wire [3:0] SAXISCCTREADY_OUT;
  wire [3:0] SAXISRQTREADY_OUT;
  wire [4:0] CFGMSGRECEIVEDTYPE_OUT;
  wire [4:0] CFGTPHSTTADDRESS_OUT;
  wire [5:0] CFGFUNCTIONPOWERSTATE_OUT;
  wire [5:0] CFGINTERRUPTMSIMMENABLE_OUT;
  wire [5:0] CFGINTERRUPTMSIVFENABLE_OUT;
  wire [5:0] CFGINTERRUPTMSIXVFENABLE_OUT;
  wire [5:0] CFGINTERRUPTMSIXVFMASK_OUT;
  wire [5:0] CFGLTSSMSTATE_OUT;
  wire [5:0] CFGTPHSTMODE_OUT;
  wire [5:0] CFGVFFLRINPROCESS_OUT;
  wire [5:0] CFGVFTPHREQUESTERENABLE_OUT;
  wire [5:0] PCIECQNPREQCOUNT_OUT;
  wire [5:0] PCIERQTAG_OUT;
  wire [5:0] PIPERX0EQLPLFFS_OUT;
  wire [5:0] PIPERX1EQLPLFFS_OUT;
  wire [5:0] PIPERX2EQLPLFFS_OUT;
  wire [5:0] PIPERX3EQLPLFFS_OUT;
  wire [5:0] PIPERX4EQLPLFFS_OUT;
  wire [5:0] PIPERX5EQLPLFFS_OUT;
  wire [5:0] PIPERX6EQLPLFFS_OUT;
  wire [5:0] PIPERX7EQLPLFFS_OUT;
  wire [5:0] PIPETX0EQDEEMPH_OUT;
  wire [5:0] PIPETX1EQDEEMPH_OUT;
  wire [5:0] PIPETX2EQDEEMPH_OUT;
  wire [5:0] PIPETX3EQDEEMPH_OUT;
  wire [5:0] PIPETX4EQDEEMPH_OUT;
  wire [5:0] PIPETX5EQDEEMPH_OUT;
  wire [5:0] PIPETX6EQDEEMPH_OUT;
  wire [5:0] PIPETX7EQDEEMPH_OUT;
  wire [71:0] MICOMPLETIONRAMWRITEDATAL_OUT;
  wire [71:0] MICOMPLETIONRAMWRITEDATAU_OUT;
  wire [74:0] MAXISRCTUSER_OUT;
  wire [7:0] CFGEXTFUNCTIONNUMBER_OUT;
  wire [7:0] CFGFCCPLH_OUT;
  wire [7:0] CFGFCNPH_OUT;
  wire [7:0] CFGFCPH_OUT;
  wire [7:0] CFGFUNCTIONSTATUS_OUT;
  wire [7:0] CFGMSGRECEIVEDDATA_OUT;
  wire [7:0] MAXISCQTKEEP_OUT;
  wire [7:0] MAXISRCTKEEP_OUT;
  wire [7:0] PLGEN3PCSRXSLIDE_OUT;
  wire [84:0] MAXISCQTUSER_OUT;
  wire [8:0] MIREPLAYRAMADDRESS_OUT;
  wire [8:0] MIREQUESTRAMREADADDRESSA_OUT;
  wire [8:0] MIREQUESTRAMREADADDRESSB_OUT;
  wire [8:0] MIREQUESTRAMWRITEADDRESSA_OUT;
  wire [8:0] MIREQUESTRAMWRITEADDRESSB_OUT;
  wire [9:0] CFGEXTREGISTERNUMBER_OUT;
  wire [9:0] MICOMPLETIONRAMREADADDRESSAL_OUT;
  wire [9:0] MICOMPLETIONRAMREADADDRESSAU_OUT;
  wire [9:0] MICOMPLETIONRAMREADADDRESSBL_OUT;
  wire [9:0] MICOMPLETIONRAMREADADDRESSBU_OUT;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSAL_OUT;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSAU_OUT;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSBL_OUT;
  wire [9:0] MICOMPLETIONRAMWRITEADDRESSBU_OUT;

  wire CFGCONFIGSPACEENABLE_IN;
  wire CFGERRCORIN_IN;
  wire CFGERRUNCORIN_IN;
  wire CFGEXTREADDATAVALID_IN;
  wire CFGHOTRESETIN_IN;
  wire CFGINPUTUPDATEREQUEST_IN;
  wire CFGINTERRUPTMSITPHPRESENT_IN;
  wire CFGINTERRUPTMSIXINT_IN;
  wire CFGLINKTRAININGENABLE_IN;
  wire CFGMCUPDATEREQUEST_IN;
  wire CFGMGMTREAD_IN;
  wire CFGMGMTTYPE1CFGREGACCESS_IN;
  wire CFGMGMTWRITE_IN;
  wire CFGMSGTRANSMIT_IN;
  wire CFGPERFUNCTIONOUTPUTREQUEST_IN;
  wire CFGPOWERSTATECHANGEACK_IN;
  wire CFGREQPMTRANSITIONL23READY_IN;
  wire CFGTPHSTTREADDATAVALID_IN;
  wire CORECLKMICOMPLETIONRAML_IN;
  wire CORECLKMICOMPLETIONRAMU_IN;
  wire CORECLKMIREPLAYRAM_IN;
  wire CORECLKMIREQUESTRAM_IN;
  wire CORECLK_IN;
  wire DRPCLK_IN;
  wire DRPEN_IN;
  wire DRPWE_IN;
  wire MGMTRESETN_IN;
  wire MGMTSTICKYRESETN_IN;
  wire PCIECQNPREQ_IN;
  wire PIPECLK_IN;
  wire PIPERESETN_IN;
  wire PIPERX0DATAVALID_IN;
  wire PIPERX0ELECIDLE_IN;
  wire PIPERX0EQDONE_IN;
  wire PIPERX0EQLPADAPTDONE_IN;
  wire PIPERX0EQLPLFFSSEL_IN;
  wire PIPERX0PHYSTATUS_IN;
  wire PIPERX0STARTBLOCK_IN;
  wire PIPERX0VALID_IN;
  wire PIPERX1DATAVALID_IN;
  wire PIPERX1ELECIDLE_IN;
  wire PIPERX1EQDONE_IN;
  wire PIPERX1EQLPADAPTDONE_IN;
  wire PIPERX1EQLPLFFSSEL_IN;
  wire PIPERX1PHYSTATUS_IN;
  wire PIPERX1STARTBLOCK_IN;
  wire PIPERX1VALID_IN;
  wire PIPERX2DATAVALID_IN;
  wire PIPERX2ELECIDLE_IN;
  wire PIPERX2EQDONE_IN;
  wire PIPERX2EQLPADAPTDONE_IN;
  wire PIPERX2EQLPLFFSSEL_IN;
  wire PIPERX2PHYSTATUS_IN;
  wire PIPERX2STARTBLOCK_IN;
  wire PIPERX2VALID_IN;
  wire PIPERX3DATAVALID_IN;
  wire PIPERX3ELECIDLE_IN;
  wire PIPERX3EQDONE_IN;
  wire PIPERX3EQLPADAPTDONE_IN;
  wire PIPERX3EQLPLFFSSEL_IN;
  wire PIPERX3PHYSTATUS_IN;
  wire PIPERX3STARTBLOCK_IN;
  wire PIPERX3VALID_IN;
  wire PIPERX4DATAVALID_IN;
  wire PIPERX4ELECIDLE_IN;
  wire PIPERX4EQDONE_IN;
  wire PIPERX4EQLPADAPTDONE_IN;
  wire PIPERX4EQLPLFFSSEL_IN;
  wire PIPERX4PHYSTATUS_IN;
  wire PIPERX4STARTBLOCK_IN;
  wire PIPERX4VALID_IN;
  wire PIPERX5DATAVALID_IN;
  wire PIPERX5ELECIDLE_IN;
  wire PIPERX5EQDONE_IN;
  wire PIPERX5EQLPADAPTDONE_IN;
  wire PIPERX5EQLPLFFSSEL_IN;
  wire PIPERX5PHYSTATUS_IN;
  wire PIPERX5STARTBLOCK_IN;
  wire PIPERX5VALID_IN;
  wire PIPERX6DATAVALID_IN;
  wire PIPERX6ELECIDLE_IN;
  wire PIPERX6EQDONE_IN;
  wire PIPERX6EQLPADAPTDONE_IN;
  wire PIPERX6EQLPLFFSSEL_IN;
  wire PIPERX6PHYSTATUS_IN;
  wire PIPERX6STARTBLOCK_IN;
  wire PIPERX6VALID_IN;
  wire PIPERX7DATAVALID_IN;
  wire PIPERX7ELECIDLE_IN;
  wire PIPERX7EQDONE_IN;
  wire PIPERX7EQLPADAPTDONE_IN;
  wire PIPERX7EQLPLFFSSEL_IN;
  wire PIPERX7PHYSTATUS_IN;
  wire PIPERX7STARTBLOCK_IN;
  wire PIPERX7VALID_IN;
  wire PIPETX0EQDONE_IN;
  wire PIPETX1EQDONE_IN;
  wire PIPETX2EQDONE_IN;
  wire PIPETX3EQDONE_IN;
  wire PIPETX4EQDONE_IN;
  wire PIPETX5EQDONE_IN;
  wire PIPETX6EQDONE_IN;
  wire PIPETX7EQDONE_IN;
  wire PLDISABLESCRAMBLER_IN;
  wire PLEQRESETEIEOSCOUNT_IN;
  wire PLGEN3PCSDISABLE_IN;
  wire RECCLK_IN;
  wire RESETN_IN;
  wire SAXISCCTLAST_IN;
  wire SAXISCCTVALID_IN;
  wire SAXISRQTLAST_IN;
  wire SAXISRQTVALID_IN;
  wire USERCLK_IN;
  wire [10:0] DRPADDR_IN;
  wire [143:0] MICOMPLETIONRAMREADDATA_IN;
  wire [143:0] MIREPLAYRAMREADDATA_IN;
  wire [143:0] MIREQUESTRAMREADDATA_IN;
  wire [15:0] CFGDEVID_IN;
  wire [15:0] CFGSUBSYSID_IN;
  wire [15:0] CFGSUBSYSVENDID_IN;
  wire [15:0] CFGVENDID_IN;
  wire [15:0] DRPDI_IN;
  wire [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET_IN;
  wire [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET_IN;
  wire [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET_IN;
  wire [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET_IN;
  wire [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET_IN;
  wire [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET_IN;
  wire [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET_IN;
  wire [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET_IN;
  wire [17:0] PIPETX0EQCOEFF_IN;
  wire [17:0] PIPETX1EQCOEFF_IN;
  wire [17:0] PIPETX2EQCOEFF_IN;
  wire [17:0] PIPETX3EQCOEFF_IN;
  wire [17:0] PIPETX4EQCOEFF_IN;
  wire [17:0] PIPETX5EQCOEFF_IN;
  wire [17:0] PIPETX6EQCOEFF_IN;
  wire [17:0] PIPETX7EQCOEFF_IN;
  wire [18:0] CFGMGMTADDR_IN;
  wire [1:0] CFGFLRDONE_IN;
  wire [1:0] CFGINTERRUPTMSITPHTYPE_IN;
  wire [1:0] CFGINTERRUPTPENDING_IN;
  wire [1:0] PIPERX0CHARISK_IN;
  wire [1:0] PIPERX0SYNCHEADER_IN;
  wire [1:0] PIPERX1CHARISK_IN;
  wire [1:0] PIPERX1SYNCHEADER_IN;
  wire [1:0] PIPERX2CHARISK_IN;
  wire [1:0] PIPERX2SYNCHEADER_IN;
  wire [1:0] PIPERX3CHARISK_IN;
  wire [1:0] PIPERX3SYNCHEADER_IN;
  wire [1:0] PIPERX4CHARISK_IN;
  wire [1:0] PIPERX4SYNCHEADER_IN;
  wire [1:0] PIPERX5CHARISK_IN;
  wire [1:0] PIPERX5SYNCHEADER_IN;
  wire [1:0] PIPERX6CHARISK_IN;
  wire [1:0] PIPERX6SYNCHEADER_IN;
  wire [1:0] PIPERX7CHARISK_IN;
  wire [1:0] PIPERX7SYNCHEADER_IN;
  wire [21:0] MAXISCQTREADY_IN;
  wire [21:0] MAXISRCTREADY_IN;
  wire [255:0] SAXISCCTDATA_IN;
  wire [255:0] SAXISRQTDATA_IN;
  wire [2:0] CFGDSFUNCTIONNUMBER_IN;
  wire [2:0] CFGFCSEL_IN;
  wire [2:0] CFGINTERRUPTMSIATTR_IN;
  wire [2:0] CFGINTERRUPTMSIFUNCTIONNUMBER_IN;
  wire [2:0] CFGMSGTRANSMITTYPE_IN;
  wire [2:0] CFGPERFUNCSTATUSCONTROL_IN;
  wire [2:0] CFGPERFUNCTIONNUMBER_IN;
  wire [2:0] PIPERX0STATUS_IN;
  wire [2:0] PIPERX1STATUS_IN;
  wire [2:0] PIPERX2STATUS_IN;
  wire [2:0] PIPERX3STATUS_IN;
  wire [2:0] PIPERX4STATUS_IN;
  wire [2:0] PIPERX5STATUS_IN;
  wire [2:0] PIPERX6STATUS_IN;
  wire [2:0] PIPERX7STATUS_IN;
  wire [31:0] CFGEXTREADDATA_IN;
  wire [31:0] CFGINTERRUPTMSIINT_IN;
  wire [31:0] CFGINTERRUPTMSIXDATA_IN;
  wire [31:0] CFGMGMTWRITEDATA_IN;
  wire [31:0] CFGMSGTRANSMITDATA_IN;
  wire [31:0] CFGTPHSTTREADDATA_IN;
  wire [31:0] PIPERX0DATA_IN;
  wire [31:0] PIPERX1DATA_IN;
  wire [31:0] PIPERX2DATA_IN;
  wire [31:0] PIPERX3DATA_IN;
  wire [31:0] PIPERX4DATA_IN;
  wire [31:0] PIPERX5DATA_IN;
  wire [31:0] PIPERX6DATA_IN;
  wire [31:0] PIPERX7DATA_IN;
  wire [32:0] SAXISCCTUSER_IN;
  wire [3:0] CFGINTERRUPTINT_IN;
  wire [3:0] CFGINTERRUPTMSISELECT_IN;
  wire [3:0] CFGMGMTBYTEENABLE_IN;
  wire [4:0] CFGDSDEVICENUMBER_IN;
  wire [59:0] SAXISRQTUSER_IN;
  wire [5:0] CFGVFFLRDONE_IN;
  wire [5:0] PIPEEQFS_IN;
  wire [5:0] PIPEEQLF_IN;
  wire [63:0] CFGDSN_IN;
  wire [63:0] CFGINTERRUPTMSIPENDINGSTATUS_IN;
  wire [63:0] CFGINTERRUPTMSIXADDRESS_IN;
  wire [7:0] CFGDSBUSNUMBER_IN;
  wire [7:0] CFGDSPORTNUMBER_IN;
  wire [7:0] CFGREVID_IN;
  wire [7:0] PLGEN3PCSRXSYNCDONE_IN;
  wire [7:0] SAXISCCTKEEP_IN;
  wire [7:0] SAXISRQTKEEP_IN;
  wire [8:0] CFGINTERRUPTMSITPHSTTAG_IN;

  wire CFGCONFIGSPACEENABLE_INDELAY;
  wire CFGERRCORIN_INDELAY;
  wire CFGERRUNCORIN_INDELAY;
  wire CFGEXTREADDATAVALID_INDELAY;
  wire CFGHOTRESETIN_INDELAY;
  wire CFGINPUTUPDATEREQUEST_INDELAY;
  wire CFGINTERRUPTMSITPHPRESENT_INDELAY;
  wire CFGINTERRUPTMSIXINT_INDELAY;
  wire CFGLINKTRAININGENABLE_INDELAY;
  wire CFGMCUPDATEREQUEST_INDELAY;
  wire CFGMGMTREAD_INDELAY;
  wire CFGMGMTTYPE1CFGREGACCESS_INDELAY;
  wire CFGMGMTWRITE_INDELAY;
  wire CFGMSGTRANSMIT_INDELAY;
  wire CFGPERFUNCTIONOUTPUTREQUEST_INDELAY;
  wire CFGPOWERSTATECHANGEACK_INDELAY;
  wire CFGREQPMTRANSITIONL23READY_INDELAY;
  wire CFGTPHSTTREADDATAVALID_INDELAY;
  wire CORECLKMICOMPLETIONRAML_INDELAY;
  wire CORECLKMICOMPLETIONRAMU_INDELAY;
  wire CORECLKMIREPLAYRAM_INDELAY;
  wire CORECLKMIREQUESTRAM_INDELAY;
  wire CORECLK_INDELAY;
  wire DRPCLK_INDELAY;
  wire DRPEN_INDELAY;
  wire DRPWE_INDELAY;
  wire MGMTRESETN_INDELAY;
  wire MGMTSTICKYRESETN_INDELAY;
  wire PCIECQNPREQ_INDELAY;
  wire PIPECLK_INDELAY;
  wire PIPERESETN_INDELAY;
  wire PIPERX0DATAVALID_INDELAY;
  wire PIPERX0ELECIDLE_INDELAY;
  wire PIPERX0EQDONE_INDELAY;
  wire PIPERX0EQLPADAPTDONE_INDELAY;
  wire PIPERX0EQLPLFFSSEL_INDELAY;
  wire PIPERX0PHYSTATUS_INDELAY;
  wire PIPERX0STARTBLOCK_INDELAY;
  wire PIPERX0VALID_INDELAY;
  wire PIPERX1DATAVALID_INDELAY;
  wire PIPERX1ELECIDLE_INDELAY;
  wire PIPERX1EQDONE_INDELAY;
  wire PIPERX1EQLPADAPTDONE_INDELAY;
  wire PIPERX1EQLPLFFSSEL_INDELAY;
  wire PIPERX1PHYSTATUS_INDELAY;
  wire PIPERX1STARTBLOCK_INDELAY;
  wire PIPERX1VALID_INDELAY;
  wire PIPERX2DATAVALID_INDELAY;
  wire PIPERX2ELECIDLE_INDELAY;
  wire PIPERX2EQDONE_INDELAY;
  wire PIPERX2EQLPADAPTDONE_INDELAY;
  wire PIPERX2EQLPLFFSSEL_INDELAY;
  wire PIPERX2PHYSTATUS_INDELAY;
  wire PIPERX2STARTBLOCK_INDELAY;
  wire PIPERX2VALID_INDELAY;
  wire PIPERX3DATAVALID_INDELAY;
  wire PIPERX3ELECIDLE_INDELAY;
  wire PIPERX3EQDONE_INDELAY;
  wire PIPERX3EQLPADAPTDONE_INDELAY;
  wire PIPERX3EQLPLFFSSEL_INDELAY;
  wire PIPERX3PHYSTATUS_INDELAY;
  wire PIPERX3STARTBLOCK_INDELAY;
  wire PIPERX3VALID_INDELAY;
  wire PIPERX4DATAVALID_INDELAY;
  wire PIPERX4ELECIDLE_INDELAY;
  wire PIPERX4EQDONE_INDELAY;
  wire PIPERX4EQLPADAPTDONE_INDELAY;
  wire PIPERX4EQLPLFFSSEL_INDELAY;
  wire PIPERX4PHYSTATUS_INDELAY;
  wire PIPERX4STARTBLOCK_INDELAY;
  wire PIPERX4VALID_INDELAY;
  wire PIPERX5DATAVALID_INDELAY;
  wire PIPERX5ELECIDLE_INDELAY;
  wire PIPERX5EQDONE_INDELAY;
  wire PIPERX5EQLPADAPTDONE_INDELAY;
  wire PIPERX5EQLPLFFSSEL_INDELAY;
  wire PIPERX5PHYSTATUS_INDELAY;
  wire PIPERX5STARTBLOCK_INDELAY;
  wire PIPERX5VALID_INDELAY;
  wire PIPERX6DATAVALID_INDELAY;
  wire PIPERX6ELECIDLE_INDELAY;
  wire PIPERX6EQDONE_INDELAY;
  wire PIPERX6EQLPADAPTDONE_INDELAY;
  wire PIPERX6EQLPLFFSSEL_INDELAY;
  wire PIPERX6PHYSTATUS_INDELAY;
  wire PIPERX6STARTBLOCK_INDELAY;
  wire PIPERX6VALID_INDELAY;
  wire PIPERX7DATAVALID_INDELAY;
  wire PIPERX7ELECIDLE_INDELAY;
  wire PIPERX7EQDONE_INDELAY;
  wire PIPERX7EQLPADAPTDONE_INDELAY;
  wire PIPERX7EQLPLFFSSEL_INDELAY;
  wire PIPERX7PHYSTATUS_INDELAY;
  wire PIPERX7STARTBLOCK_INDELAY;
  wire PIPERX7VALID_INDELAY;
  wire PIPETX0EQDONE_INDELAY;
  wire PIPETX1EQDONE_INDELAY;
  wire PIPETX2EQDONE_INDELAY;
  wire PIPETX3EQDONE_INDELAY;
  wire PIPETX4EQDONE_INDELAY;
  wire PIPETX5EQDONE_INDELAY;
  wire PIPETX6EQDONE_INDELAY;
  wire PIPETX7EQDONE_INDELAY;
  wire PLDISABLESCRAMBLER_INDELAY;
  wire PLEQRESETEIEOSCOUNT_INDELAY;
  wire PLGEN3PCSDISABLE_INDELAY;
  wire RECCLK_INDELAY;
  wire RESETN_INDELAY;
  wire SAXISCCTLAST_INDELAY;
  wire SAXISCCTVALID_INDELAY;
  wire SAXISRQTLAST_INDELAY;
  wire SAXISRQTVALID_INDELAY;
  wire USERCLK_INDELAY;
  wire [10:0] DRPADDR_INDELAY;
  wire [143:0] MICOMPLETIONRAMREADDATA_INDELAY;
  wire [143:0] MIREPLAYRAMREADDATA_INDELAY;
  wire [143:0] MIREQUESTRAMREADDATA_INDELAY;
  wire [15:0] CFGDEVID_INDELAY;
  wire [15:0] CFGSUBSYSID_INDELAY;
  wire [15:0] CFGSUBSYSVENDID_INDELAY;
  wire [15:0] CFGVENDID_INDELAY;
  wire [15:0] DRPDI_INDELAY;
  wire [17:0] PIPERX0EQLPNEWTXCOEFFORPRESET_INDELAY;
  wire [17:0] PIPERX1EQLPNEWTXCOEFFORPRESET_INDELAY;
  wire [17:0] PIPERX2EQLPNEWTXCOEFFORPRESET_INDELAY;
  wire [17:0] PIPERX3EQLPNEWTXCOEFFORPRESET_INDELAY;
  wire [17:0] PIPERX4EQLPNEWTXCOEFFORPRESET_INDELAY;
  wire [17:0] PIPERX5EQLPNEWTXCOEFFORPRESET_INDELAY;
  wire [17:0] PIPERX6EQLPNEWTXCOEFFORPRESET_INDELAY;
  wire [17:0] PIPERX7EQLPNEWTXCOEFFORPRESET_INDELAY;
  wire [17:0] PIPETX0EQCOEFF_INDELAY;
  wire [17:0] PIPETX1EQCOEFF_INDELAY;
  wire [17:0] PIPETX2EQCOEFF_INDELAY;
  wire [17:0] PIPETX3EQCOEFF_INDELAY;
  wire [17:0] PIPETX4EQCOEFF_INDELAY;
  wire [17:0] PIPETX5EQCOEFF_INDELAY;
  wire [17:0] PIPETX6EQCOEFF_INDELAY;
  wire [17:0] PIPETX7EQCOEFF_INDELAY;
  wire [18:0] CFGMGMTADDR_INDELAY;
  wire [1:0] CFGFLRDONE_INDELAY;
  wire [1:0] CFGINTERRUPTMSITPHTYPE_INDELAY;
  wire [1:0] CFGINTERRUPTPENDING_INDELAY;
  wire [1:0] PIPERX0CHARISK_INDELAY;
  wire [1:0] PIPERX0SYNCHEADER_INDELAY;
  wire [1:0] PIPERX1CHARISK_INDELAY;
  wire [1:0] PIPERX1SYNCHEADER_INDELAY;
  wire [1:0] PIPERX2CHARISK_INDELAY;
  wire [1:0] PIPERX2SYNCHEADER_INDELAY;
  wire [1:0] PIPERX3CHARISK_INDELAY;
  wire [1:0] PIPERX3SYNCHEADER_INDELAY;
  wire [1:0] PIPERX4CHARISK_INDELAY;
  wire [1:0] PIPERX4SYNCHEADER_INDELAY;
  wire [1:0] PIPERX5CHARISK_INDELAY;
  wire [1:0] PIPERX5SYNCHEADER_INDELAY;
  wire [1:0] PIPERX6CHARISK_INDELAY;
  wire [1:0] PIPERX6SYNCHEADER_INDELAY;
  wire [1:0] PIPERX7CHARISK_INDELAY;
  wire [1:0] PIPERX7SYNCHEADER_INDELAY;
  wire [21:0] MAXISCQTREADY_INDELAY;
  wire [21:0] MAXISRCTREADY_INDELAY;
  wire [255:0] SAXISCCTDATA_INDELAY;
  wire [255:0] SAXISRQTDATA_INDELAY;
  wire [2:0] CFGDSFUNCTIONNUMBER_INDELAY;
  wire [2:0] CFGFCSEL_INDELAY;
  wire [2:0] CFGINTERRUPTMSIATTR_INDELAY;
  wire [2:0] CFGINTERRUPTMSIFUNCTIONNUMBER_INDELAY;
  wire [2:0] CFGMSGTRANSMITTYPE_INDELAY;
  wire [2:0] CFGPERFUNCSTATUSCONTROL_INDELAY;
  wire [2:0] CFGPERFUNCTIONNUMBER_INDELAY;
  wire [2:0] PIPERX0STATUS_INDELAY;
  wire [2:0] PIPERX1STATUS_INDELAY;
  wire [2:0] PIPERX2STATUS_INDELAY;
  wire [2:0] PIPERX3STATUS_INDELAY;
  wire [2:0] PIPERX4STATUS_INDELAY;
  wire [2:0] PIPERX5STATUS_INDELAY;
  wire [2:0] PIPERX6STATUS_INDELAY;
  wire [2:0] PIPERX7STATUS_INDELAY;
  wire [31:0] CFGEXTREADDATA_INDELAY;
  wire [31:0] CFGINTERRUPTMSIINT_INDELAY;
  wire [31:0] CFGINTERRUPTMSIXDATA_INDELAY;
  wire [31:0] CFGMGMTWRITEDATA_INDELAY;
  wire [31:0] CFGMSGTRANSMITDATA_INDELAY;
  wire [31:0] CFGTPHSTTREADDATA_INDELAY;
  wire [31:0] PIPERX0DATA_INDELAY;
  wire [31:0] PIPERX1DATA_INDELAY;
  wire [31:0] PIPERX2DATA_INDELAY;
  wire [31:0] PIPERX3DATA_INDELAY;
  wire [31:0] PIPERX4DATA_INDELAY;
  wire [31:0] PIPERX5DATA_INDELAY;
  wire [31:0] PIPERX6DATA_INDELAY;
  wire [31:0] PIPERX7DATA_INDELAY;
  wire [32:0] SAXISCCTUSER_INDELAY;
  wire [3:0] CFGINTERRUPTINT_INDELAY;
  wire [3:0] CFGINTERRUPTMSISELECT_INDELAY;
  wire [3:0] CFGMGMTBYTEENABLE_INDELAY;
  wire [4:0] CFGDSDEVICENUMBER_INDELAY;
  wire [59:0] SAXISRQTUSER_INDELAY;
  wire [5:0] CFGVFFLRDONE_INDELAY;
  wire [5:0] PIPEEQFS_INDELAY;
  wire [5:0] PIPEEQLF_INDELAY;
  wire [63:0] CFGDSN_INDELAY;
  wire [63:0] CFGINTERRUPTMSIPENDINGSTATUS_INDELAY;
  wire [63:0] CFGINTERRUPTMSIXADDRESS_INDELAY;
  wire [7:0] CFGDSBUSNUMBER_INDELAY;
  wire [7:0] CFGDSPORTNUMBER_INDELAY;
  wire [7:0] CFGREVID_INDELAY;
  wire [7:0] PLGEN3PCSRXSYNCDONE_INDELAY;
  wire [7:0] SAXISCCTKEEP_INDELAY;
  wire [7:0] SAXISRQTKEEP_INDELAY;
  wire [8:0] CFGINTERRUPTMSITPHSTTAG_INDELAY;

  initial begin
    case (ARI_CAP_ENABLE)
      "FALSE" : ARI_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : ARI_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute ARI_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", ARI_CAP_ENABLE);
        $finish;
      end
    endcase

    case (AXISTEN_IF_CC_ALIGNMENT_MODE)
      "FALSE" : AXISTEN_IF_CC_ALIGNMENT_MODE_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_CC_ALIGNMENT_MODE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_CC_ALIGNMENT_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_CC_ALIGNMENT_MODE);
        $finish;
      end
    endcase

    case (AXISTEN_IF_CC_PARITY_CHK)
      "TRUE" : AXISTEN_IF_CC_PARITY_CHK_BINARY = 1'b1;
      "FALSE" : AXISTEN_IF_CC_PARITY_CHK_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_CC_PARITY_CHK on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", AXISTEN_IF_CC_PARITY_CHK);
        $finish;
      end
    endcase

    case (AXISTEN_IF_CQ_ALIGNMENT_MODE)
      "FALSE" : AXISTEN_IF_CQ_ALIGNMENT_MODE_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_CQ_ALIGNMENT_MODE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_CQ_ALIGNMENT_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_CQ_ALIGNMENT_MODE);
        $finish;
      end
    endcase

    case (AXISTEN_IF_ENABLE_CLIENT_TAG)
      "FALSE" : AXISTEN_IF_ENABLE_CLIENT_TAG_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_ENABLE_CLIENT_TAG_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_ENABLE_CLIENT_TAG on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_ENABLE_CLIENT_TAG);
        $finish;
      end
    endcase

    case (AXISTEN_IF_ENABLE_RX_MSG_INTFC)
      "FALSE" : AXISTEN_IF_ENABLE_RX_MSG_INTFC_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_ENABLE_RX_MSG_INTFC_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_ENABLE_RX_MSG_INTFC on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_ENABLE_RX_MSG_INTFC);
        $finish;
      end
    endcase

    case (AXISTEN_IF_RC_ALIGNMENT_MODE)
      "FALSE" : AXISTEN_IF_RC_ALIGNMENT_MODE_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_RC_ALIGNMENT_MODE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_RC_ALIGNMENT_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_RC_ALIGNMENT_MODE);
        $finish;
      end
    endcase

    case (AXISTEN_IF_RC_STRADDLE)
      "FALSE" : AXISTEN_IF_RC_STRADDLE_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_RC_STRADDLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_RC_STRADDLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_RC_STRADDLE);
        $finish;
      end
    endcase

    case (AXISTEN_IF_RQ_ALIGNMENT_MODE)
      "FALSE" : AXISTEN_IF_RQ_ALIGNMENT_MODE_BINARY = 1'b0;
      "TRUE" : AXISTEN_IF_RQ_ALIGNMENT_MODE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_RQ_ALIGNMENT_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", AXISTEN_IF_RQ_ALIGNMENT_MODE);
        $finish;
      end
    endcase

    case (AXISTEN_IF_RQ_PARITY_CHK)
      "TRUE" : AXISTEN_IF_RQ_PARITY_CHK_BINARY = 1'b1;
      "FALSE" : AXISTEN_IF_RQ_PARITY_CHK_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute AXISTEN_IF_RQ_PARITY_CHK on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", AXISTEN_IF_RQ_PARITY_CHK);
        $finish;
      end
    endcase

    case (CRM_CORE_CLK_FREQ_500)
      "TRUE" : CRM_CORE_CLK_FREQ_500_BINARY = 1'b1;
      "FALSE" : CRM_CORE_CLK_FREQ_500_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute CRM_CORE_CLK_FREQ_500 on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", CRM_CORE_CLK_FREQ_500);
        $finish;
      end
    endcase

    case (GEN3_PCS_RX_ELECIDLE_INTERNAL)
      "TRUE" : GEN3_PCS_RX_ELECIDLE_INTERNAL_BINARY = 1'b1;
      "FALSE" : GEN3_PCS_RX_ELECIDLE_INTERNAL_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute GEN3_PCS_RX_ELECIDLE_INTERNAL on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", GEN3_PCS_RX_ELECIDLE_INTERNAL);
        $finish;
      end
    endcase

    case (LL_ACK_TIMEOUT_EN)
      "FALSE" : LL_ACK_TIMEOUT_EN_BINARY = 1'b0;
      "TRUE" : LL_ACK_TIMEOUT_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_ACK_TIMEOUT_EN on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_ACK_TIMEOUT_EN);
        $finish;
      end
    endcase

    case (LL_CPL_FC_UPDATE_TIMER_OVERRIDE)
      "FALSE" : LL_CPL_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b0;
      "TRUE" : LL_CPL_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_CPL_FC_UPDATE_TIMER_OVERRIDE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_CPL_FC_UPDATE_TIMER_OVERRIDE);
        $finish;
      end
    endcase

    case (LL_FC_UPDATE_TIMER_OVERRIDE)
      "FALSE" : LL_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b0;
      "TRUE" : LL_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_FC_UPDATE_TIMER_OVERRIDE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_FC_UPDATE_TIMER_OVERRIDE);
        $finish;
      end
    endcase

    case (LL_NP_FC_UPDATE_TIMER_OVERRIDE)
      "FALSE" : LL_NP_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b0;
      "TRUE" : LL_NP_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_NP_FC_UPDATE_TIMER_OVERRIDE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_NP_FC_UPDATE_TIMER_OVERRIDE);
        $finish;
      end
    endcase

    case (LL_P_FC_UPDATE_TIMER_OVERRIDE)
      "FALSE" : LL_P_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b0;
      "TRUE" : LL_P_FC_UPDATE_TIMER_OVERRIDE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_P_FC_UPDATE_TIMER_OVERRIDE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_P_FC_UPDATE_TIMER_OVERRIDE);
        $finish;
      end
    endcase

    case (LL_REPLAY_TIMEOUT_EN)
      "FALSE" : LL_REPLAY_TIMEOUT_EN_BINARY = 1'b0;
      "TRUE" : LL_REPLAY_TIMEOUT_EN_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LL_REPLAY_TIMEOUT_EN on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LL_REPLAY_TIMEOUT_EN);
        $finish;
      end
    endcase

    case (LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE)
      "FALSE" : LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_BINARY = 1'b0;
      "TRUE" : LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE);
        $finish;
      end
    endcase

    case (LTR_TX_MESSAGE_ON_LTR_ENABLE)
      "FALSE" : LTR_TX_MESSAGE_ON_LTR_ENABLE_BINARY = 1'b0;
      "TRUE" : LTR_TX_MESSAGE_ON_LTR_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute LTR_TX_MESSAGE_ON_LTR_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", LTR_TX_MESSAGE_ON_LTR_ENABLE);
        $finish;
      end
    endcase

    case (PF0_AER_CAP_ECRC_CHECK_CAPABLE)
      "FALSE" : PF0_AER_CAP_ECRC_CHECK_CAPABLE_BINARY = 1'b0;
      "TRUE" : PF0_AER_CAP_ECRC_CHECK_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_AER_CAP_ECRC_CHECK_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_AER_CAP_ECRC_CHECK_CAPABLE);
        $finish;
      end
    endcase

    case (PF0_AER_CAP_ECRC_GEN_CAPABLE)
      "FALSE" : PF0_AER_CAP_ECRC_GEN_CAPABLE_BINARY = 1'b0;
      "TRUE" : PF0_AER_CAP_ECRC_GEN_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_AER_CAP_ECRC_GEN_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_AER_CAP_ECRC_GEN_CAPABLE);
        $finish;
      end
    endcase

    case (PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT)
      "TRUE" : PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT);
        $finish;
      end
    endcase

    case (PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT)
      "TRUE" : PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT);
        $finish;
      end
    endcase

    case (PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT)
      "TRUE" : PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT);
        $finish;
      end
    endcase

    case (PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE)
      "TRUE" : PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE);
        $finish;
      end
    endcase

    case (PF0_DEV_CAP2_LTR_SUPPORT)
      "TRUE" : PF0_DEV_CAP2_LTR_SUPPORT_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP2_LTR_SUPPORT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_LTR_SUPPORT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP2_LTR_SUPPORT);
        $finish;
      end
    endcase

    case (PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT)
      "FALSE" : PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_BINARY = 1'b0;
      "TRUE" : PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT);
        $finish;
      end
    endcase

    case (PF0_DEV_CAP_EXT_TAG_SUPPORTED)
      "TRUE" : PF0_DEV_CAP_EXT_TAG_SUPPORTED_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP_EXT_TAG_SUPPORTED_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP_EXT_TAG_SUPPORTED on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP_EXT_TAG_SUPPORTED);
        $finish;
      end
    endcase

    case (PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE)
      "TRUE" : PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_BINARY = 1'b1;
      "FALSE" : PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE);
        $finish;
      end
    endcase

    case (PF0_DPA_CAP_SUB_STATE_CONTROL_EN)
      "TRUE" : PF0_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY = 1'b1;
      "FALSE" : PF0_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_DPA_CAP_SUB_STATE_CONTROL_EN on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_DPA_CAP_SUB_STATE_CONTROL_EN);
        $finish;
      end
    endcase

    case (PF0_EXPANSION_ROM_ENABLE)
      "FALSE" : PF0_EXPANSION_ROM_ENABLE_BINARY = 1'b0;
      "TRUE" : PF0_EXPANSION_ROM_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_EXPANSION_ROM_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_EXPANSION_ROM_ENABLE);
        $finish;
      end
    endcase

    case (PF0_LINK_STATUS_SLOT_CLOCK_CONFIG)
      "TRUE" : PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_BINARY = 1'b1;
      "FALSE" : PF0_LINK_STATUS_SLOT_CLOCK_CONFIG_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_LINK_STATUS_SLOT_CLOCK_CONFIG on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_LINK_STATUS_SLOT_CLOCK_CONFIG);
        $finish;
      end
    endcase

    case (PF0_PB_CAP_SYSTEM_ALLOCATED)
      "FALSE" : PF0_PB_CAP_SYSTEM_ALLOCATED_BINARY = 1'b0;
      "TRUE" : PF0_PB_CAP_SYSTEM_ALLOCATED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PB_CAP_SYSTEM_ALLOCATED on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_PB_CAP_SYSTEM_ALLOCATED);
        $finish;
      end
    endcase

    case (PF0_PM_CAP_PMESUPPORT_D0)
      "TRUE" : PF0_PM_CAP_PMESUPPORT_D0_BINARY = 1'b1;
      "FALSE" : PF0_PM_CAP_PMESUPPORT_D0_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PM_CAP_PMESUPPORT_D0 on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_PM_CAP_PMESUPPORT_D0);
        $finish;
      end
    endcase

    case (PF0_PM_CAP_PMESUPPORT_D1)
      "TRUE" : PF0_PM_CAP_PMESUPPORT_D1_BINARY = 1'b1;
      "FALSE" : PF0_PM_CAP_PMESUPPORT_D1_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PM_CAP_PMESUPPORT_D1 on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_PM_CAP_PMESUPPORT_D1);
        $finish;
      end
    endcase

    case (PF0_PM_CAP_PMESUPPORT_D3HOT)
      "TRUE" : PF0_PM_CAP_PMESUPPORT_D3HOT_BINARY = 1'b1;
      "FALSE" : PF0_PM_CAP_PMESUPPORT_D3HOT_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PM_CAP_PMESUPPORT_D3HOT on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_PM_CAP_PMESUPPORT_D3HOT);
        $finish;
      end
    endcase

    case (PF0_PM_CAP_SUPP_D1_STATE)
      "TRUE" : PF0_PM_CAP_SUPP_D1_STATE_BINARY = 1'b1;
      "FALSE" : PF0_PM_CAP_SUPP_D1_STATE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PM_CAP_SUPP_D1_STATE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_PM_CAP_SUPP_D1_STATE);
        $finish;
      end
    endcase

    case (PF0_PM_CSR_NOSOFTRESET)
      "TRUE" : PF0_PM_CSR_NOSOFTRESET_BINARY = 1'b1;
      "FALSE" : PF0_PM_CSR_NOSOFTRESET_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_PM_CSR_NOSOFTRESET on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_PM_CSR_NOSOFTRESET);
        $finish;
      end
    endcase

    case (PF0_RBAR_CAP_ENABLE)
      "FALSE" : PF0_RBAR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : PF0_RBAR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_RBAR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_RBAR_CAP_ENABLE);
        $finish;
      end
    endcase

    case (PF0_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : PF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : PF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_TPHR_CAP_DEV_SPECIFIC_MODE);
        $finish;
      end
    endcase

    case (PF0_TPHR_CAP_ENABLE)
      "FALSE" : PF0_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : PF0_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF0_TPHR_CAP_ENABLE);
        $finish;
      end
    endcase

    case (PF0_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : PF0_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : PF0_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF0_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF0_TPHR_CAP_INT_VEC_MODE);
        $finish;
      end
    endcase

    case (PF1_AER_CAP_ECRC_CHECK_CAPABLE)
      "FALSE" : PF1_AER_CAP_ECRC_CHECK_CAPABLE_BINARY = 1'b0;
      "TRUE" : PF1_AER_CAP_ECRC_CHECK_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_AER_CAP_ECRC_CHECK_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_AER_CAP_ECRC_CHECK_CAPABLE);
        $finish;
      end
    endcase

    case (PF1_AER_CAP_ECRC_GEN_CAPABLE)
      "FALSE" : PF1_AER_CAP_ECRC_GEN_CAPABLE_BINARY = 1'b0;
      "TRUE" : PF1_AER_CAP_ECRC_GEN_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_AER_CAP_ECRC_GEN_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_AER_CAP_ECRC_GEN_CAPABLE);
        $finish;
      end
    endcase

    case (PF1_DPA_CAP_SUB_STATE_CONTROL_EN)
      "TRUE" : PF1_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY = 1'b1;
      "FALSE" : PF1_DPA_CAP_SUB_STATE_CONTROL_EN_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_DPA_CAP_SUB_STATE_CONTROL_EN on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF1_DPA_CAP_SUB_STATE_CONTROL_EN);
        $finish;
      end
    endcase

    case (PF1_EXPANSION_ROM_ENABLE)
      "FALSE" : PF1_EXPANSION_ROM_ENABLE_BINARY = 1'b0;
      "TRUE" : PF1_EXPANSION_ROM_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_EXPANSION_ROM_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_EXPANSION_ROM_ENABLE);
        $finish;
      end
    endcase

    case (PF1_PB_CAP_SYSTEM_ALLOCATED)
      "FALSE" : PF1_PB_CAP_SYSTEM_ALLOCATED_BINARY = 1'b0;
      "TRUE" : PF1_PB_CAP_SYSTEM_ALLOCATED_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_PB_CAP_SYSTEM_ALLOCATED on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_PB_CAP_SYSTEM_ALLOCATED);
        $finish;
      end
    endcase

    case (PF1_RBAR_CAP_ENABLE)
      "FALSE" : PF1_RBAR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : PF1_RBAR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_RBAR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_RBAR_CAP_ENABLE);
        $finish;
      end
    endcase

    case (PF1_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : PF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : PF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF1_TPHR_CAP_DEV_SPECIFIC_MODE);
        $finish;
      end
    endcase

    case (PF1_TPHR_CAP_ENABLE)
      "FALSE" : PF1_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : PF1_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PF1_TPHR_CAP_ENABLE);
        $finish;
      end
    endcase

    case (PF1_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : PF1_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : PF1_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PF1_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PF1_TPHR_CAP_INT_VEC_MODE);
        $finish;
      end
    endcase

    case (PL_DISABLE_EI_INFER_IN_L0)
      "FALSE" : PL_DISABLE_EI_INFER_IN_L0_BINARY = 1'b0;
      "TRUE" : PL_DISABLE_EI_INFER_IN_L0_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_DISABLE_EI_INFER_IN_L0 on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_DISABLE_EI_INFER_IN_L0);
        $finish;
      end
    endcase

    case (PL_DISABLE_GEN3_DC_BALANCE)
      "FALSE" : PL_DISABLE_GEN3_DC_BALANCE_BINARY = 1'b0;
      "TRUE" : PL_DISABLE_GEN3_DC_BALANCE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_DISABLE_GEN3_DC_BALANCE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_DISABLE_GEN3_DC_BALANCE);
        $finish;
      end
    endcase

    case (PL_DISABLE_SCRAMBLING)
      "FALSE" : PL_DISABLE_SCRAMBLING_BINARY = 1'b0;
      "TRUE" : PL_DISABLE_SCRAMBLING_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_DISABLE_SCRAMBLING on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_DISABLE_SCRAMBLING);
        $finish;
      end
    endcase

    case (PL_DISABLE_UPCONFIG_CAPABLE)
      "FALSE" : PL_DISABLE_UPCONFIG_CAPABLE_BINARY = 1'b0;
      "TRUE" : PL_DISABLE_UPCONFIG_CAPABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_DISABLE_UPCONFIG_CAPABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_DISABLE_UPCONFIG_CAPABLE);
        $finish;
      end
    endcase

    case (PL_EQ_ADAPT_DISABLE_COEFF_CHECK)
      "FALSE" : PL_EQ_ADAPT_DISABLE_COEFF_CHECK_BINARY = 1'b0;
      "TRUE" : PL_EQ_ADAPT_DISABLE_COEFF_CHECK_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_EQ_ADAPT_DISABLE_COEFF_CHECK on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_EQ_ADAPT_DISABLE_COEFF_CHECK);
        $finish;
      end
    endcase

    case (PL_EQ_ADAPT_DISABLE_PRESET_CHECK)
      "FALSE" : PL_EQ_ADAPT_DISABLE_PRESET_CHECK_BINARY = 1'b0;
      "TRUE" : PL_EQ_ADAPT_DISABLE_PRESET_CHECK_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_EQ_ADAPT_DISABLE_PRESET_CHECK on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_EQ_ADAPT_DISABLE_PRESET_CHECK);
        $finish;
      end
    endcase

    case (PL_EQ_BYPASS_PHASE23)
      "FALSE" : PL_EQ_BYPASS_PHASE23_BINARY = 1'b0;
      "TRUE" : PL_EQ_BYPASS_PHASE23_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_EQ_BYPASS_PHASE23 on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_EQ_BYPASS_PHASE23);
        $finish;
      end
    endcase

    case (PL_EQ_SHORT_ADAPT_PHASE)
      "FALSE" : PL_EQ_SHORT_ADAPT_PHASE_BINARY = 1'b0;
      "TRUE" : PL_EQ_SHORT_ADAPT_PHASE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_EQ_SHORT_ADAPT_PHASE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_EQ_SHORT_ADAPT_PHASE);
        $finish;
      end
    endcase

    case (PL_SIM_FAST_LINK_TRAINING)
      "FALSE" : PL_SIM_FAST_LINK_TRAINING_BINARY = 1'b0;
      "TRUE" : PL_SIM_FAST_LINK_TRAINING_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_SIM_FAST_LINK_TRAINING on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", PL_SIM_FAST_LINK_TRAINING);
        $finish;
      end
    endcase

    case (PL_UPSTREAM_FACING)
      "TRUE" : PL_UPSTREAM_FACING_BINARY = 1'b1;
      "FALSE" : PL_UPSTREAM_FACING_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PL_UPSTREAM_FACING on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PL_UPSTREAM_FACING);
        $finish;
      end
    endcase

    case (PM_ENABLE_SLOT_POWER_CAPTURE)
      "TRUE" : PM_ENABLE_SLOT_POWER_CAPTURE_BINARY = 1'b1;
      "FALSE" : PM_ENABLE_SLOT_POWER_CAPTURE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute PM_ENABLE_SLOT_POWER_CAPTURE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", PM_ENABLE_SLOT_POWER_CAPTURE);
        $finish;
      end
    endcase

    case (SIM_VERSION)
      "1.0" : SIM_VERSION_BINARY = 0;
      "1.1" : SIM_VERSION_BINARY = 0;
      "1.2" : SIM_VERSION_BINARY = 0;
      "1.3" : SIM_VERSION_BINARY = 0;
      "2.0" : SIM_VERSION_BINARY = 0;
      "3.0" : SIM_VERSION_BINARY = 0;
      "4.0" : SIM_VERSION_BINARY = 0;
      default : begin
        $display("Attribute Syntax Error : The Attribute SIM_VERSION on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are 1.0, 1.1, 1.2, 1.3, 2.0, 3.0, or 4.0.", SIM_VERSION);
        $finish;
      end
    endcase

    case (SRIOV_CAP_ENABLE)
      "FALSE" : SRIOV_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : SRIOV_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute SRIOV_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", SRIOV_CAP_ENABLE);
        $finish;
      end
    endcase

    case (TL_ENABLE_MESSAGE_RID_CHECK_ENABLE)
      "TRUE" : TL_ENABLE_MESSAGE_RID_CHECK_ENABLE_BINARY = 1'b1;
      "FALSE" : TL_ENABLE_MESSAGE_RID_CHECK_ENABLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_ENABLE_MESSAGE_RID_CHECK_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", TL_ENABLE_MESSAGE_RID_CHECK_ENABLE);
        $finish;
      end
    endcase

    case (TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE)
      "FALSE" : TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_BINARY = 1'b0;
      "TRUE" : TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE);
        $finish;
      end
    endcase

    case (TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE)
      "FALSE" : TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE_BINARY = 1'b0;
      "TRUE" : TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE);
        $finish;
      end
    endcase

    case (TL_LEGACY_MODE_ENABLE)
      "FALSE" : TL_LEGACY_MODE_ENABLE_BINARY = 1'b0;
      "TRUE" : TL_LEGACY_MODE_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_LEGACY_MODE_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TL_LEGACY_MODE_ENABLE);
        $finish;
      end
    endcase

    case (TL_PF_ENABLE_REG)
      "FALSE" : TL_PF_ENABLE_REG_BINARY = 1'b0;
      "TRUE" : TL_PF_ENABLE_REG_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_PF_ENABLE_REG on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", TL_PF_ENABLE_REG);
        $finish;
      end
    endcase

    case (TL_TAG_MGMT_ENABLE)
      "TRUE" : TL_TAG_MGMT_ENABLE_BINARY = 1'b1;
      "FALSE" : TL_TAG_MGMT_ENABLE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute TL_TAG_MGMT_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", TL_TAG_MGMT_ENABLE);
        $finish;
      end
    endcase

    case (VF0_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF0_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF0_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF0_TPHR_CAP_DEV_SPECIFIC_MODE);
        $finish;
      end
    endcase

    case (VF0_TPHR_CAP_ENABLE)
      "FALSE" : VF0_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF0_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF0_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF0_TPHR_CAP_ENABLE);
        $finish;
      end
    endcase

    case (VF0_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF0_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF0_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF0_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF0_TPHR_CAP_INT_VEC_MODE);
        $finish;
      end
    endcase

    case (VF1_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF1_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF1_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF1_TPHR_CAP_DEV_SPECIFIC_MODE);
        $finish;
      end
    endcase

    case (VF1_TPHR_CAP_ENABLE)
      "FALSE" : VF1_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF1_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF1_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF1_TPHR_CAP_ENABLE);
        $finish;
      end
    endcase

    case (VF1_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF1_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF1_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF1_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF1_TPHR_CAP_INT_VEC_MODE);
        $finish;
      end
    endcase

    case (VF2_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF2_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF2_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF2_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF2_TPHR_CAP_DEV_SPECIFIC_MODE);
        $finish;
      end
    endcase

    case (VF2_TPHR_CAP_ENABLE)
      "FALSE" : VF2_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF2_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF2_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF2_TPHR_CAP_ENABLE);
        $finish;
      end
    endcase

    case (VF2_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF2_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF2_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF2_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF2_TPHR_CAP_INT_VEC_MODE);
        $finish;
      end
    endcase

    case (VF3_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF3_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF3_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF3_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF3_TPHR_CAP_DEV_SPECIFIC_MODE);
        $finish;
      end
    endcase

    case (VF3_TPHR_CAP_ENABLE)
      "FALSE" : VF3_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF3_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF3_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF3_TPHR_CAP_ENABLE);
        $finish;
      end
    endcase

    case (VF3_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF3_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF3_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF3_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF3_TPHR_CAP_INT_VEC_MODE);
        $finish;
      end
    endcase

    case (VF4_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF4_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF4_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF4_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF4_TPHR_CAP_DEV_SPECIFIC_MODE);
        $finish;
      end
    endcase

    case (VF4_TPHR_CAP_ENABLE)
      "FALSE" : VF4_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF4_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF4_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF4_TPHR_CAP_ENABLE);
        $finish;
      end
    endcase

    case (VF4_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF4_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF4_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF4_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF4_TPHR_CAP_INT_VEC_MODE);
        $finish;
      end
    endcase

    case (VF5_TPHR_CAP_DEV_SPECIFIC_MODE)
      "TRUE" : VF5_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b1;
      "FALSE" : VF5_TPHR_CAP_DEV_SPECIFIC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF5_TPHR_CAP_DEV_SPECIFIC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF5_TPHR_CAP_DEV_SPECIFIC_MODE);
        $finish;
      end
    endcase

    case (VF5_TPHR_CAP_ENABLE)
      "FALSE" : VF5_TPHR_CAP_ENABLE_BINARY = 1'b0;
      "TRUE" : VF5_TPHR_CAP_ENABLE_BINARY = 1'b1;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF5_TPHR_CAP_ENABLE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are FALSE, or TRUE.", VF5_TPHR_CAP_ENABLE);
        $finish;
      end
    endcase

    case (VF5_TPHR_CAP_INT_VEC_MODE)
      "TRUE" : VF5_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b1;
      "FALSE" : VF5_TPHR_CAP_INT_VEC_MODE_BINARY = 1'b0;
      default : begin
        $display("Attribute Syntax Error : The Attribute VF5_TPHR_CAP_INT_VEC_MODE on X_PCIE_3_0 instance %m is set to %s.  Legal values for this attribute are TRUE, or FALSE.", VF5_TPHR_CAP_INT_VEC_MODE);
        $finish;
      end
    endcase

    if ((LL_ACK_TIMEOUT_FUNC >= 0) && (LL_ACK_TIMEOUT_FUNC <= 3))
      LL_ACK_TIMEOUT_FUNC_BINARY = LL_ACK_TIMEOUT_FUNC;
    else begin
      $display("Attribute Syntax Error : The Attribute LL_ACK_TIMEOUT_FUNC on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", LL_ACK_TIMEOUT_FUNC);
      $finish;
    end

    if ((LL_REPLAY_TIMEOUT_FUNC >= 0) && (LL_REPLAY_TIMEOUT_FUNC <= 3))
      LL_REPLAY_TIMEOUT_FUNC_BINARY = LL_REPLAY_TIMEOUT_FUNC;
    else begin
      $display("Attribute Syntax Error : The Attribute LL_REPLAY_TIMEOUT_FUNC on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", LL_REPLAY_TIMEOUT_FUNC);
      $finish;
    end

    if ((PF0_DEV_CAP_ENDPOINT_L0S_LATENCY >= 0) && (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY <= 7))
      PF0_DEV_CAP_ENDPOINT_L0S_LATENCY_BINARY = PF0_DEV_CAP_ENDPOINT_L0S_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP_ENDPOINT_L0S_LATENCY on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_DEV_CAP_ENDPOINT_L0S_LATENCY);
      $finish;
    end

    if ((PF0_DEV_CAP_ENDPOINT_L1_LATENCY >= 0) && (PF0_DEV_CAP_ENDPOINT_L1_LATENCY <= 7))
      PF0_DEV_CAP_ENDPOINT_L1_LATENCY_BINARY = PF0_DEV_CAP_ENDPOINT_L1_LATENCY;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_DEV_CAP_ENDPOINT_L1_LATENCY on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_DEV_CAP_ENDPOINT_L1_LATENCY);
      $finish;
    end

    if ((PF0_LINK_CAP_ASPM_SUPPORT >= 0) && (PF0_LINK_CAP_ASPM_SUPPORT <= 3))
      PF0_LINK_CAP_ASPM_SUPPORT_BINARY = PF0_LINK_CAP_ASPM_SUPPORT;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_ASPM_SUPPORT on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 3.", PF0_LINK_CAP_ASPM_SUPPORT);
      $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1);
      $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2);
      $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3);
      $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1);
      $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2);
      $finish;
    end

    if ((PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 >= 0) && (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 <= 7))
      PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3_BINARY = PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3);
      $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1);
      $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2);
      $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3);
      $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1);
      $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2);
      $finish;
    end

    if ((PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 >= 0) && (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 <= 7))
      PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3_BINARY = PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3);
      $finish;
    end

    if ((PF0_MSIX_CAP_PBA_BIR >= 0) && (PF0_MSIX_CAP_PBA_BIR <= 7))
      PF0_MSIX_CAP_PBA_BIR_BINARY = PF0_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_MSIX_CAP_PBA_BIR);
      $finish;
    end

    if ((PF0_MSIX_CAP_TABLE_BIR >= 0) && (PF0_MSIX_CAP_TABLE_BIR <= 7))
      PF0_MSIX_CAP_TABLE_BIR_BINARY = PF0_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_MSIX_CAP_TABLE_BIR);
      $finish;
    end

    if ((PF0_MSI_CAP_MULTIMSGCAP >= 0) && (PF0_MSI_CAP_MULTIMSGCAP <= 7))
      PF0_MSI_CAP_MULTIMSGCAP_BINARY = PF0_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute PF0_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF0_MSI_CAP_MULTIMSGCAP);
      $finish;
    end

    if ((PF1_MSIX_CAP_PBA_BIR >= 0) && (PF1_MSIX_CAP_PBA_BIR <= 7))
      PF1_MSIX_CAP_PBA_BIR_BINARY = PF1_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute PF1_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF1_MSIX_CAP_PBA_BIR);
      $finish;
    end

    if ((PF1_MSIX_CAP_TABLE_BIR >= 0) && (PF1_MSIX_CAP_TABLE_BIR <= 7))
      PF1_MSIX_CAP_TABLE_BIR_BINARY = PF1_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute PF1_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF1_MSIX_CAP_TABLE_BIR);
      $finish;
    end

    if ((PF1_MSI_CAP_MULTIMSGCAP >= 0) && (PF1_MSI_CAP_MULTIMSGCAP <= 7))
      PF1_MSI_CAP_MULTIMSGCAP_BINARY = PF1_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute PF1_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", PF1_MSI_CAP_MULTIMSGCAP);
      $finish;
    end

    if ((PL_N_FTS_COMCLK_GEN1 >= 0) && (PL_N_FTS_COMCLK_GEN1 <= 255))
      PL_N_FTS_COMCLK_GEN1_BINARY = PL_N_FTS_COMCLK_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_COMCLK_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_COMCLK_GEN1);
      $finish;
    end

    if ((PL_N_FTS_COMCLK_GEN2 >= 0) && (PL_N_FTS_COMCLK_GEN2 <= 255))
      PL_N_FTS_COMCLK_GEN2_BINARY = PL_N_FTS_COMCLK_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_COMCLK_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_COMCLK_GEN2);
      $finish;
    end

    if ((PL_N_FTS_COMCLK_GEN3 >= 0) && (PL_N_FTS_COMCLK_GEN3 <= 255))
      PL_N_FTS_COMCLK_GEN3_BINARY = PL_N_FTS_COMCLK_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_COMCLK_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_COMCLK_GEN3);
      $finish;
    end

    if ((PL_N_FTS_GEN1 >= 0) && (PL_N_FTS_GEN1 <= 255))
      PL_N_FTS_GEN1_BINARY = PL_N_FTS_GEN1;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_GEN1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_GEN1);
      $finish;
    end

    if ((PL_N_FTS_GEN2 >= 0) && (PL_N_FTS_GEN2 <= 255))
      PL_N_FTS_GEN2_BINARY = PL_N_FTS_GEN2;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_GEN2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_GEN2);
      $finish;
    end

    if ((PL_N_FTS_GEN3 >= 0) && (PL_N_FTS_GEN3 <= 255))
      PL_N_FTS_GEN3_BINARY = PL_N_FTS_GEN3;
    else begin
      $display("Attribute Syntax Error : The Attribute PL_N_FTS_GEN3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 255.", PL_N_FTS_GEN3);
      $finish;
    end

    if ((SPARE_BIT0 >= 0) && (SPARE_BIT0 <= 1))
      SPARE_BIT0_BINARY = SPARE_BIT0;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT0 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT0);
      $finish;
    end

    if ((SPARE_BIT1 >= 0) && (SPARE_BIT1 <= 1))
      SPARE_BIT1_BINARY = SPARE_BIT1;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT1 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT1);
      $finish;
    end

    if ((SPARE_BIT2 >= 0) && (SPARE_BIT2 <= 1))
      SPARE_BIT2_BINARY = SPARE_BIT2;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT2 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT2);
      $finish;
    end

    if ((SPARE_BIT3 >= 0) && (SPARE_BIT3 <= 1))
      SPARE_BIT3_BINARY = SPARE_BIT3;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT3 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT3);
      $finish;
    end

    if ((SPARE_BIT4 >= 0) && (SPARE_BIT4 <= 1))
      SPARE_BIT4_BINARY = SPARE_BIT4;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT4 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT4);
      $finish;
    end

    if ((SPARE_BIT5 >= 0) && (SPARE_BIT5 <= 1))
      SPARE_BIT5_BINARY = SPARE_BIT5;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT5 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT5);
      $finish;
    end

    if ((SPARE_BIT6 >= 0) && (SPARE_BIT6 <= 1))
      SPARE_BIT6_BINARY = SPARE_BIT6;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT6 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT6);
      $finish;
    end

    if ((SPARE_BIT7 >= 0) && (SPARE_BIT7 <= 1))
      SPARE_BIT7_BINARY = SPARE_BIT7;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT7 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT7);
      $finish;
    end

    if ((SPARE_BIT8 >= 0) && (SPARE_BIT8 <= 1))
      SPARE_BIT8_BINARY = SPARE_BIT8;
    else begin
      $display("Attribute Syntax Error : The Attribute SPARE_BIT8 on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 1.", SPARE_BIT8);
      $finish;
    end

    if ((VF0_MSIX_CAP_PBA_BIR >= 0) && (VF0_MSIX_CAP_PBA_BIR <= 7))
      VF0_MSIX_CAP_PBA_BIR_BINARY = VF0_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF0_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF0_MSIX_CAP_PBA_BIR);
      $finish;
    end

    if ((VF0_MSIX_CAP_TABLE_BIR >= 0) && (VF0_MSIX_CAP_TABLE_BIR <= 7))
      VF0_MSIX_CAP_TABLE_BIR_BINARY = VF0_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF0_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF0_MSIX_CAP_TABLE_BIR);
      $finish;
    end

    if ((VF0_MSI_CAP_MULTIMSGCAP >= 0) && (VF0_MSI_CAP_MULTIMSGCAP <= 7))
      VF0_MSI_CAP_MULTIMSGCAP_BINARY = VF0_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF0_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF0_MSI_CAP_MULTIMSGCAP);
      $finish;
    end

    if ((VF1_MSIX_CAP_PBA_BIR >= 0) && (VF1_MSIX_CAP_PBA_BIR <= 7))
      VF1_MSIX_CAP_PBA_BIR_BINARY = VF1_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF1_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF1_MSIX_CAP_PBA_BIR);
      $finish;
    end

    if ((VF1_MSIX_CAP_TABLE_BIR >= 0) && (VF1_MSIX_CAP_TABLE_BIR <= 7))
      VF1_MSIX_CAP_TABLE_BIR_BINARY = VF1_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF1_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF1_MSIX_CAP_TABLE_BIR);
      $finish;
    end

    if ((VF1_MSI_CAP_MULTIMSGCAP >= 0) && (VF1_MSI_CAP_MULTIMSGCAP <= 7))
      VF1_MSI_CAP_MULTIMSGCAP_BINARY = VF1_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF1_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF1_MSI_CAP_MULTIMSGCAP);
      $finish;
    end

    if ((VF2_MSIX_CAP_PBA_BIR >= 0) && (VF2_MSIX_CAP_PBA_BIR <= 7))
      VF2_MSIX_CAP_PBA_BIR_BINARY = VF2_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF2_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF2_MSIX_CAP_PBA_BIR);
      $finish;
    end

    if ((VF2_MSIX_CAP_TABLE_BIR >= 0) && (VF2_MSIX_CAP_TABLE_BIR <= 7))
      VF2_MSIX_CAP_TABLE_BIR_BINARY = VF2_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF2_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF2_MSIX_CAP_TABLE_BIR);
      $finish;
    end

    if ((VF2_MSI_CAP_MULTIMSGCAP >= 0) && (VF2_MSI_CAP_MULTIMSGCAP <= 7))
      VF2_MSI_CAP_MULTIMSGCAP_BINARY = VF2_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF2_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF2_MSI_CAP_MULTIMSGCAP);
      $finish;
    end

    if ((VF3_MSIX_CAP_PBA_BIR >= 0) && (VF3_MSIX_CAP_PBA_BIR <= 7))
      VF3_MSIX_CAP_PBA_BIR_BINARY = VF3_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF3_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF3_MSIX_CAP_PBA_BIR);
      $finish;
    end

    if ((VF3_MSIX_CAP_TABLE_BIR >= 0) && (VF3_MSIX_CAP_TABLE_BIR <= 7))
      VF3_MSIX_CAP_TABLE_BIR_BINARY = VF3_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF3_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF3_MSIX_CAP_TABLE_BIR);
      $finish;
    end

    if ((VF3_MSI_CAP_MULTIMSGCAP >= 0) && (VF3_MSI_CAP_MULTIMSGCAP <= 7))
      VF3_MSI_CAP_MULTIMSGCAP_BINARY = VF3_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF3_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF3_MSI_CAP_MULTIMSGCAP);
      $finish;
    end

    if ((VF4_MSIX_CAP_PBA_BIR >= 0) && (VF4_MSIX_CAP_PBA_BIR <= 7))
      VF4_MSIX_CAP_PBA_BIR_BINARY = VF4_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF4_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF4_MSIX_CAP_PBA_BIR);
      $finish;
    end

    if ((VF4_MSIX_CAP_TABLE_BIR >= 0) && (VF4_MSIX_CAP_TABLE_BIR <= 7))
      VF4_MSIX_CAP_TABLE_BIR_BINARY = VF4_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF4_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF4_MSIX_CAP_TABLE_BIR);
      $finish;
    end

    if ((VF4_MSI_CAP_MULTIMSGCAP >= 0) && (VF4_MSI_CAP_MULTIMSGCAP <= 7))
      VF4_MSI_CAP_MULTIMSGCAP_BINARY = VF4_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF4_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF4_MSI_CAP_MULTIMSGCAP);
      $finish;
    end

    if ((VF5_MSIX_CAP_PBA_BIR >= 0) && (VF5_MSIX_CAP_PBA_BIR <= 7))
      VF5_MSIX_CAP_PBA_BIR_BINARY = VF5_MSIX_CAP_PBA_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF5_MSIX_CAP_PBA_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF5_MSIX_CAP_PBA_BIR);
      $finish;
    end

    if ((VF5_MSIX_CAP_TABLE_BIR >= 0) && (VF5_MSIX_CAP_TABLE_BIR <= 7))
      VF5_MSIX_CAP_TABLE_BIR_BINARY = VF5_MSIX_CAP_TABLE_BIR;
    else begin
      $display("Attribute Syntax Error : The Attribute VF5_MSIX_CAP_TABLE_BIR on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF5_MSIX_CAP_TABLE_BIR);
      $finish;
    end

    if ((VF5_MSI_CAP_MULTIMSGCAP >= 0) && (VF5_MSI_CAP_MULTIMSGCAP <= 7))
      VF5_MSI_CAP_MULTIMSGCAP_BINARY = VF5_MSI_CAP_MULTIMSGCAP;
    else begin
      $display("Attribute Syntax Error : The Attribute VF5_MSI_CAP_MULTIMSGCAP on X_PCIE_3_0 instance %m is set to %d.  Legal values for this attribute are  0 to 7.", VF5_MSI_CAP_MULTIMSGCAP);
      $finish;
    end

  end

  buf B_CFGCURRENTSPEED0 (CFGCURRENTSPEED[0], CFGCURRENTSPEED_OUT[0]);
  buf B_CFGCURRENTSPEED1 (CFGCURRENTSPEED[1], CFGCURRENTSPEED_OUT[1]);
  buf B_CFGCURRENTSPEED2 (CFGCURRENTSPEED[2], CFGCURRENTSPEED_OUT[2]);
  buf B_CFGDPASUBSTATECHANGE0 (CFGDPASUBSTATECHANGE[0], CFGDPASUBSTATECHANGE_OUT[0]);
  buf B_CFGDPASUBSTATECHANGE1 (CFGDPASUBSTATECHANGE[1], CFGDPASUBSTATECHANGE_OUT[1]);
  buf B_CFGERRCOROUT (CFGERRCOROUT, CFGERRCOROUT_OUT);
  buf B_CFGERRFATALOUT (CFGERRFATALOUT, CFGERRFATALOUT_OUT);
  buf B_CFGERRNONFATALOUT (CFGERRNONFATALOUT, CFGERRNONFATALOUT_OUT);
  buf B_CFGEXTFUNCTIONNUMBER0 (CFGEXTFUNCTIONNUMBER[0], CFGEXTFUNCTIONNUMBER_OUT[0]);
  buf B_CFGEXTFUNCTIONNUMBER1 (CFGEXTFUNCTIONNUMBER[1], CFGEXTFUNCTIONNUMBER_OUT[1]);
  buf B_CFGEXTFUNCTIONNUMBER2 (CFGEXTFUNCTIONNUMBER[2], CFGEXTFUNCTIONNUMBER_OUT[2]);
  buf B_CFGEXTFUNCTIONNUMBER3 (CFGEXTFUNCTIONNUMBER[3], CFGEXTFUNCTIONNUMBER_OUT[3]);
  buf B_CFGEXTFUNCTIONNUMBER4 (CFGEXTFUNCTIONNUMBER[4], CFGEXTFUNCTIONNUMBER_OUT[4]);
  buf B_CFGEXTFUNCTIONNUMBER5 (CFGEXTFUNCTIONNUMBER[5], CFGEXTFUNCTIONNUMBER_OUT[5]);
  buf B_CFGEXTFUNCTIONNUMBER6 (CFGEXTFUNCTIONNUMBER[6], CFGEXTFUNCTIONNUMBER_OUT[6]);
  buf B_CFGEXTFUNCTIONNUMBER7 (CFGEXTFUNCTIONNUMBER[7], CFGEXTFUNCTIONNUMBER_OUT[7]);
  buf B_CFGEXTREADRECEIVED (CFGEXTREADRECEIVED, CFGEXTREADRECEIVED_OUT);
  buf B_CFGEXTREGISTERNUMBER0 (CFGEXTREGISTERNUMBER[0], CFGEXTREGISTERNUMBER_OUT[0]);
  buf B_CFGEXTREGISTERNUMBER1 (CFGEXTREGISTERNUMBER[1], CFGEXTREGISTERNUMBER_OUT[1]);
  buf B_CFGEXTREGISTERNUMBER2 (CFGEXTREGISTERNUMBER[2], CFGEXTREGISTERNUMBER_OUT[2]);
  buf B_CFGEXTREGISTERNUMBER3 (CFGEXTREGISTERNUMBER[3], CFGEXTREGISTERNUMBER_OUT[3]);
  buf B_CFGEXTREGISTERNUMBER4 (CFGEXTREGISTERNUMBER[4], CFGEXTREGISTERNUMBER_OUT[4]);
  buf B_CFGEXTREGISTERNUMBER5 (CFGEXTREGISTERNUMBER[5], CFGEXTREGISTERNUMBER_OUT[5]);
  buf B_CFGEXTREGISTERNUMBER6 (CFGEXTREGISTERNUMBER[6], CFGEXTREGISTERNUMBER_OUT[6]);
  buf B_CFGEXTREGISTERNUMBER7 (CFGEXTREGISTERNUMBER[7], CFGEXTREGISTERNUMBER_OUT[7]);
  buf B_CFGEXTREGISTERNUMBER8 (CFGEXTREGISTERNUMBER[8], CFGEXTREGISTERNUMBER_OUT[8]);
  buf B_CFGEXTREGISTERNUMBER9 (CFGEXTREGISTERNUMBER[9], CFGEXTREGISTERNUMBER_OUT[9]);
  buf B_CFGEXTWRITEBYTEENABLE0 (CFGEXTWRITEBYTEENABLE[0], CFGEXTWRITEBYTEENABLE_OUT[0]);
  buf B_CFGEXTWRITEBYTEENABLE1 (CFGEXTWRITEBYTEENABLE[1], CFGEXTWRITEBYTEENABLE_OUT[1]);
  buf B_CFGEXTWRITEBYTEENABLE2 (CFGEXTWRITEBYTEENABLE[2], CFGEXTWRITEBYTEENABLE_OUT[2]);
  buf B_CFGEXTWRITEBYTEENABLE3 (CFGEXTWRITEBYTEENABLE[3], CFGEXTWRITEBYTEENABLE_OUT[3]);
  buf B_CFGEXTWRITEDATA0 (CFGEXTWRITEDATA[0], CFGEXTWRITEDATA_OUT[0]);
  buf B_CFGEXTWRITEDATA1 (CFGEXTWRITEDATA[1], CFGEXTWRITEDATA_OUT[1]);
  buf B_CFGEXTWRITEDATA10 (CFGEXTWRITEDATA[10], CFGEXTWRITEDATA_OUT[10]);
  buf B_CFGEXTWRITEDATA11 (CFGEXTWRITEDATA[11], CFGEXTWRITEDATA_OUT[11]);
  buf B_CFGEXTWRITEDATA12 (CFGEXTWRITEDATA[12], CFGEXTWRITEDATA_OUT[12]);
  buf B_CFGEXTWRITEDATA13 (CFGEXTWRITEDATA[13], CFGEXTWRITEDATA_OUT[13]);
  buf B_CFGEXTWRITEDATA14 (CFGEXTWRITEDATA[14], CFGEXTWRITEDATA_OUT[14]);
  buf B_CFGEXTWRITEDATA15 (CFGEXTWRITEDATA[15], CFGEXTWRITEDATA_OUT[15]);
  buf B_CFGEXTWRITEDATA16 (CFGEXTWRITEDATA[16], CFGEXTWRITEDATA_OUT[16]);
  buf B_CFGEXTWRITEDATA17 (CFGEXTWRITEDATA[17], CFGEXTWRITEDATA_OUT[17]);
  buf B_CFGEXTWRITEDATA18 (CFGEXTWRITEDATA[18], CFGEXTWRITEDATA_OUT[18]);
  buf B_CFGEXTWRITEDATA19 (CFGEXTWRITEDATA[19], CFGEXTWRITEDATA_OUT[19]);
  buf B_CFGEXTWRITEDATA2 (CFGEXTWRITEDATA[2], CFGEXTWRITEDATA_OUT[2]);
  buf B_CFGEXTWRITEDATA20 (CFGEXTWRITEDATA[20], CFGEXTWRITEDATA_OUT[20]);
  buf B_CFGEXTWRITEDATA21 (CFGEXTWRITEDATA[21], CFGEXTWRITEDATA_OUT[21]);
  buf B_CFGEXTWRITEDATA22 (CFGEXTWRITEDATA[22], CFGEXTWRITEDATA_OUT[22]);
  buf B_CFGEXTWRITEDATA23 (CFGEXTWRITEDATA[23], CFGEXTWRITEDATA_OUT[23]);
  buf B_CFGEXTWRITEDATA24 (CFGEXTWRITEDATA[24], CFGEXTWRITEDATA_OUT[24]);
  buf B_CFGEXTWRITEDATA25 (CFGEXTWRITEDATA[25], CFGEXTWRITEDATA_OUT[25]);
  buf B_CFGEXTWRITEDATA26 (CFGEXTWRITEDATA[26], CFGEXTWRITEDATA_OUT[26]);
  buf B_CFGEXTWRITEDATA27 (CFGEXTWRITEDATA[27], CFGEXTWRITEDATA_OUT[27]);
  buf B_CFGEXTWRITEDATA28 (CFGEXTWRITEDATA[28], CFGEXTWRITEDATA_OUT[28]);
  buf B_CFGEXTWRITEDATA29 (CFGEXTWRITEDATA[29], CFGEXTWRITEDATA_OUT[29]);
  buf B_CFGEXTWRITEDATA3 (CFGEXTWRITEDATA[3], CFGEXTWRITEDATA_OUT[3]);
  buf B_CFGEXTWRITEDATA30 (CFGEXTWRITEDATA[30], CFGEXTWRITEDATA_OUT[30]);
  buf B_CFGEXTWRITEDATA31 (CFGEXTWRITEDATA[31], CFGEXTWRITEDATA_OUT[31]);
  buf B_CFGEXTWRITEDATA4 (CFGEXTWRITEDATA[4], CFGEXTWRITEDATA_OUT[4]);
  buf B_CFGEXTWRITEDATA5 (CFGEXTWRITEDATA[5], CFGEXTWRITEDATA_OUT[5]);
  buf B_CFGEXTWRITEDATA6 (CFGEXTWRITEDATA[6], CFGEXTWRITEDATA_OUT[6]);
  buf B_CFGEXTWRITEDATA7 (CFGEXTWRITEDATA[7], CFGEXTWRITEDATA_OUT[7]);
  buf B_CFGEXTWRITEDATA8 (CFGEXTWRITEDATA[8], CFGEXTWRITEDATA_OUT[8]);
  buf B_CFGEXTWRITEDATA9 (CFGEXTWRITEDATA[9], CFGEXTWRITEDATA_OUT[9]);
  buf B_CFGEXTWRITERECEIVED (CFGEXTWRITERECEIVED, CFGEXTWRITERECEIVED_OUT);
  buf B_CFGFCCPLD0 (CFGFCCPLD[0], CFGFCCPLD_OUT[0]);
  buf B_CFGFCCPLD1 (CFGFCCPLD[1], CFGFCCPLD_OUT[1]);
  buf B_CFGFCCPLD10 (CFGFCCPLD[10], CFGFCCPLD_OUT[10]);
  buf B_CFGFCCPLD11 (CFGFCCPLD[11], CFGFCCPLD_OUT[11]);
  buf B_CFGFCCPLD2 (CFGFCCPLD[2], CFGFCCPLD_OUT[2]);
  buf B_CFGFCCPLD3 (CFGFCCPLD[3], CFGFCCPLD_OUT[3]);
  buf B_CFGFCCPLD4 (CFGFCCPLD[4], CFGFCCPLD_OUT[4]);
  buf B_CFGFCCPLD5 (CFGFCCPLD[5], CFGFCCPLD_OUT[5]);
  buf B_CFGFCCPLD6 (CFGFCCPLD[6], CFGFCCPLD_OUT[6]);
  buf B_CFGFCCPLD7 (CFGFCCPLD[7], CFGFCCPLD_OUT[7]);
  buf B_CFGFCCPLD8 (CFGFCCPLD[8], CFGFCCPLD_OUT[8]);
  buf B_CFGFCCPLD9 (CFGFCCPLD[9], CFGFCCPLD_OUT[9]);
  buf B_CFGFCCPLH0 (CFGFCCPLH[0], CFGFCCPLH_OUT[0]);
  buf B_CFGFCCPLH1 (CFGFCCPLH[1], CFGFCCPLH_OUT[1]);
  buf B_CFGFCCPLH2 (CFGFCCPLH[2], CFGFCCPLH_OUT[2]);
  buf B_CFGFCCPLH3 (CFGFCCPLH[3], CFGFCCPLH_OUT[3]);
  buf B_CFGFCCPLH4 (CFGFCCPLH[4], CFGFCCPLH_OUT[4]);
  buf B_CFGFCCPLH5 (CFGFCCPLH[5], CFGFCCPLH_OUT[5]);
  buf B_CFGFCCPLH6 (CFGFCCPLH[6], CFGFCCPLH_OUT[6]);
  buf B_CFGFCCPLH7 (CFGFCCPLH[7], CFGFCCPLH_OUT[7]);
  buf B_CFGFCNPD0 (CFGFCNPD[0], CFGFCNPD_OUT[0]);
  buf B_CFGFCNPD1 (CFGFCNPD[1], CFGFCNPD_OUT[1]);
  buf B_CFGFCNPD10 (CFGFCNPD[10], CFGFCNPD_OUT[10]);
  buf B_CFGFCNPD11 (CFGFCNPD[11], CFGFCNPD_OUT[11]);
  buf B_CFGFCNPD2 (CFGFCNPD[2], CFGFCNPD_OUT[2]);
  buf B_CFGFCNPD3 (CFGFCNPD[3], CFGFCNPD_OUT[3]);
  buf B_CFGFCNPD4 (CFGFCNPD[4], CFGFCNPD_OUT[4]);
  buf B_CFGFCNPD5 (CFGFCNPD[5], CFGFCNPD_OUT[5]);
  buf B_CFGFCNPD6 (CFGFCNPD[6], CFGFCNPD_OUT[6]);
  buf B_CFGFCNPD7 (CFGFCNPD[7], CFGFCNPD_OUT[7]);
  buf B_CFGFCNPD8 (CFGFCNPD[8], CFGFCNPD_OUT[8]);
  buf B_CFGFCNPD9 (CFGFCNPD[9], CFGFCNPD_OUT[9]);
  buf B_CFGFCNPH0 (CFGFCNPH[0], CFGFCNPH_OUT[0]);
  buf B_CFGFCNPH1 (CFGFCNPH[1], CFGFCNPH_OUT[1]);
  buf B_CFGFCNPH2 (CFGFCNPH[2], CFGFCNPH_OUT[2]);
  buf B_CFGFCNPH3 (CFGFCNPH[3], CFGFCNPH_OUT[3]);
  buf B_CFGFCNPH4 (CFGFCNPH[4], CFGFCNPH_OUT[4]);
  buf B_CFGFCNPH5 (CFGFCNPH[5], CFGFCNPH_OUT[5]);
  buf B_CFGFCNPH6 (CFGFCNPH[6], CFGFCNPH_OUT[6]);
  buf B_CFGFCNPH7 (CFGFCNPH[7], CFGFCNPH_OUT[7]);
  buf B_CFGFCPD0 (CFGFCPD[0], CFGFCPD_OUT[0]);
  buf B_CFGFCPD1 (CFGFCPD[1], CFGFCPD_OUT[1]);
  buf B_CFGFCPD10 (CFGFCPD[10], CFGFCPD_OUT[10]);
  buf B_CFGFCPD11 (CFGFCPD[11], CFGFCPD_OUT[11]);
  buf B_CFGFCPD2 (CFGFCPD[2], CFGFCPD_OUT[2]);
  buf B_CFGFCPD3 (CFGFCPD[3], CFGFCPD_OUT[3]);
  buf B_CFGFCPD4 (CFGFCPD[4], CFGFCPD_OUT[4]);
  buf B_CFGFCPD5 (CFGFCPD[5], CFGFCPD_OUT[5]);
  buf B_CFGFCPD6 (CFGFCPD[6], CFGFCPD_OUT[6]);
  buf B_CFGFCPD7 (CFGFCPD[7], CFGFCPD_OUT[7]);
  buf B_CFGFCPD8 (CFGFCPD[8], CFGFCPD_OUT[8]);
  buf B_CFGFCPD9 (CFGFCPD[9], CFGFCPD_OUT[9]);
  buf B_CFGFCPH0 (CFGFCPH[0], CFGFCPH_OUT[0]);
  buf B_CFGFCPH1 (CFGFCPH[1], CFGFCPH_OUT[1]);
  buf B_CFGFCPH2 (CFGFCPH[2], CFGFCPH_OUT[2]);
  buf B_CFGFCPH3 (CFGFCPH[3], CFGFCPH_OUT[3]);
  buf B_CFGFCPH4 (CFGFCPH[4], CFGFCPH_OUT[4]);
  buf B_CFGFCPH5 (CFGFCPH[5], CFGFCPH_OUT[5]);
  buf B_CFGFCPH6 (CFGFCPH[6], CFGFCPH_OUT[6]);
  buf B_CFGFCPH7 (CFGFCPH[7], CFGFCPH_OUT[7]);
  buf B_CFGFLRINPROCESS0 (CFGFLRINPROCESS[0], CFGFLRINPROCESS_OUT[0]);
  buf B_CFGFLRINPROCESS1 (CFGFLRINPROCESS[1], CFGFLRINPROCESS_OUT[1]);
  buf B_CFGFUNCTIONPOWERSTATE0 (CFGFUNCTIONPOWERSTATE[0], CFGFUNCTIONPOWERSTATE_OUT[0]);
  buf B_CFGFUNCTIONPOWERSTATE1 (CFGFUNCTIONPOWERSTATE[1], CFGFUNCTIONPOWERSTATE_OUT[1]);
  buf B_CFGFUNCTIONPOWERSTATE2 (CFGFUNCTIONPOWERSTATE[2], CFGFUNCTIONPOWERSTATE_OUT[2]);
  buf B_CFGFUNCTIONPOWERSTATE3 (CFGFUNCTIONPOWERSTATE[3], CFGFUNCTIONPOWERSTATE_OUT[3]);
  buf B_CFGFUNCTIONPOWERSTATE4 (CFGFUNCTIONPOWERSTATE[4], CFGFUNCTIONPOWERSTATE_OUT[4]);
  buf B_CFGFUNCTIONPOWERSTATE5 (CFGFUNCTIONPOWERSTATE[5], CFGFUNCTIONPOWERSTATE_OUT[5]);
  buf B_CFGFUNCTIONSTATUS0 (CFGFUNCTIONSTATUS[0], CFGFUNCTIONSTATUS_OUT[0]);
  buf B_CFGFUNCTIONSTATUS1 (CFGFUNCTIONSTATUS[1], CFGFUNCTIONSTATUS_OUT[1]);
  buf B_CFGFUNCTIONSTATUS2 (CFGFUNCTIONSTATUS[2], CFGFUNCTIONSTATUS_OUT[2]);
  buf B_CFGFUNCTIONSTATUS3 (CFGFUNCTIONSTATUS[3], CFGFUNCTIONSTATUS_OUT[3]);
  buf B_CFGFUNCTIONSTATUS4 (CFGFUNCTIONSTATUS[4], CFGFUNCTIONSTATUS_OUT[4]);
  buf B_CFGFUNCTIONSTATUS5 (CFGFUNCTIONSTATUS[5], CFGFUNCTIONSTATUS_OUT[5]);
  buf B_CFGFUNCTIONSTATUS6 (CFGFUNCTIONSTATUS[6], CFGFUNCTIONSTATUS_OUT[6]);
  buf B_CFGFUNCTIONSTATUS7 (CFGFUNCTIONSTATUS[7], CFGFUNCTIONSTATUS_OUT[7]);
  buf B_CFGHOTRESETOUT (CFGHOTRESETOUT, CFGHOTRESETOUT_OUT);
  buf B_CFGINPUTUPDATEDONE (CFGINPUTUPDATEDONE, CFGINPUTUPDATEDONE_OUT);
  buf B_CFGINTERRUPTAOUTPUT (CFGINTERRUPTAOUTPUT, CFGINTERRUPTAOUTPUT_OUT);
  buf B_CFGINTERRUPTBOUTPUT (CFGINTERRUPTBOUTPUT, CFGINTERRUPTBOUTPUT_OUT);
  buf B_CFGINTERRUPTCOUTPUT (CFGINTERRUPTCOUTPUT, CFGINTERRUPTCOUTPUT_OUT);
  buf B_CFGINTERRUPTDOUTPUT (CFGINTERRUPTDOUTPUT, CFGINTERRUPTDOUTPUT_OUT);
  buf B_CFGINTERRUPTMSIDATA0 (CFGINTERRUPTMSIDATA[0], CFGINTERRUPTMSIDATA_OUT[0]);
  buf B_CFGINTERRUPTMSIDATA1 (CFGINTERRUPTMSIDATA[1], CFGINTERRUPTMSIDATA_OUT[1]);
  buf B_CFGINTERRUPTMSIDATA10 (CFGINTERRUPTMSIDATA[10], CFGINTERRUPTMSIDATA_OUT[10]);
  buf B_CFGINTERRUPTMSIDATA11 (CFGINTERRUPTMSIDATA[11], CFGINTERRUPTMSIDATA_OUT[11]);
  buf B_CFGINTERRUPTMSIDATA12 (CFGINTERRUPTMSIDATA[12], CFGINTERRUPTMSIDATA_OUT[12]);
  buf B_CFGINTERRUPTMSIDATA13 (CFGINTERRUPTMSIDATA[13], CFGINTERRUPTMSIDATA_OUT[13]);
  buf B_CFGINTERRUPTMSIDATA14 (CFGINTERRUPTMSIDATA[14], CFGINTERRUPTMSIDATA_OUT[14]);
  buf B_CFGINTERRUPTMSIDATA15 (CFGINTERRUPTMSIDATA[15], CFGINTERRUPTMSIDATA_OUT[15]);
  buf B_CFGINTERRUPTMSIDATA16 (CFGINTERRUPTMSIDATA[16], CFGINTERRUPTMSIDATA_OUT[16]);
  buf B_CFGINTERRUPTMSIDATA17 (CFGINTERRUPTMSIDATA[17], CFGINTERRUPTMSIDATA_OUT[17]);
  buf B_CFGINTERRUPTMSIDATA18 (CFGINTERRUPTMSIDATA[18], CFGINTERRUPTMSIDATA_OUT[18]);
  buf B_CFGINTERRUPTMSIDATA19 (CFGINTERRUPTMSIDATA[19], CFGINTERRUPTMSIDATA_OUT[19]);
  buf B_CFGINTERRUPTMSIDATA2 (CFGINTERRUPTMSIDATA[2], CFGINTERRUPTMSIDATA_OUT[2]);
  buf B_CFGINTERRUPTMSIDATA20 (CFGINTERRUPTMSIDATA[20], CFGINTERRUPTMSIDATA_OUT[20]);
  buf B_CFGINTERRUPTMSIDATA21 (CFGINTERRUPTMSIDATA[21], CFGINTERRUPTMSIDATA_OUT[21]);
  buf B_CFGINTERRUPTMSIDATA22 (CFGINTERRUPTMSIDATA[22], CFGINTERRUPTMSIDATA_OUT[22]);
  buf B_CFGINTERRUPTMSIDATA23 (CFGINTERRUPTMSIDATA[23], CFGINTERRUPTMSIDATA_OUT[23]);
  buf B_CFGINTERRUPTMSIDATA24 (CFGINTERRUPTMSIDATA[24], CFGINTERRUPTMSIDATA_OUT[24]);
  buf B_CFGINTERRUPTMSIDATA25 (CFGINTERRUPTMSIDATA[25], CFGINTERRUPTMSIDATA_OUT[25]);
  buf B_CFGINTERRUPTMSIDATA26 (CFGINTERRUPTMSIDATA[26], CFGINTERRUPTMSIDATA_OUT[26]);
  buf B_CFGINTERRUPTMSIDATA27 (CFGINTERRUPTMSIDATA[27], CFGINTERRUPTMSIDATA_OUT[27]);
  buf B_CFGINTERRUPTMSIDATA28 (CFGINTERRUPTMSIDATA[28], CFGINTERRUPTMSIDATA_OUT[28]);
  buf B_CFGINTERRUPTMSIDATA29 (CFGINTERRUPTMSIDATA[29], CFGINTERRUPTMSIDATA_OUT[29]);
  buf B_CFGINTERRUPTMSIDATA3 (CFGINTERRUPTMSIDATA[3], CFGINTERRUPTMSIDATA_OUT[3]);
  buf B_CFGINTERRUPTMSIDATA30 (CFGINTERRUPTMSIDATA[30], CFGINTERRUPTMSIDATA_OUT[30]);
  buf B_CFGINTERRUPTMSIDATA31 (CFGINTERRUPTMSIDATA[31], CFGINTERRUPTMSIDATA_OUT[31]);
  buf B_CFGINTERRUPTMSIDATA4 (CFGINTERRUPTMSIDATA[4], CFGINTERRUPTMSIDATA_OUT[4]);
  buf B_CFGINTERRUPTMSIDATA5 (CFGINTERRUPTMSIDATA[5], CFGINTERRUPTMSIDATA_OUT[5]);
  buf B_CFGINTERRUPTMSIDATA6 (CFGINTERRUPTMSIDATA[6], CFGINTERRUPTMSIDATA_OUT[6]);
  buf B_CFGINTERRUPTMSIDATA7 (CFGINTERRUPTMSIDATA[7], CFGINTERRUPTMSIDATA_OUT[7]);
  buf B_CFGINTERRUPTMSIDATA8 (CFGINTERRUPTMSIDATA[8], CFGINTERRUPTMSIDATA_OUT[8]);
  buf B_CFGINTERRUPTMSIDATA9 (CFGINTERRUPTMSIDATA[9], CFGINTERRUPTMSIDATA_OUT[9]);
  buf B_CFGINTERRUPTMSIENABLE0 (CFGINTERRUPTMSIENABLE[0], CFGINTERRUPTMSIENABLE_OUT[0]);
  buf B_CFGINTERRUPTMSIENABLE1 (CFGINTERRUPTMSIENABLE[1], CFGINTERRUPTMSIENABLE_OUT[1]);
  buf B_CFGINTERRUPTMSIFAIL (CFGINTERRUPTMSIFAIL, CFGINTERRUPTMSIFAIL_OUT);
  buf B_CFGINTERRUPTMSIMASKUPDATE (CFGINTERRUPTMSIMASKUPDATE, CFGINTERRUPTMSIMASKUPDATE_OUT);
  buf B_CFGINTERRUPTMSIMMENABLE0 (CFGINTERRUPTMSIMMENABLE[0], CFGINTERRUPTMSIMMENABLE_OUT[0]);
  buf B_CFGINTERRUPTMSIMMENABLE1 (CFGINTERRUPTMSIMMENABLE[1], CFGINTERRUPTMSIMMENABLE_OUT[1]);
  buf B_CFGINTERRUPTMSIMMENABLE2 (CFGINTERRUPTMSIMMENABLE[2], CFGINTERRUPTMSIMMENABLE_OUT[2]);
  buf B_CFGINTERRUPTMSIMMENABLE3 (CFGINTERRUPTMSIMMENABLE[3], CFGINTERRUPTMSIMMENABLE_OUT[3]);
  buf B_CFGINTERRUPTMSIMMENABLE4 (CFGINTERRUPTMSIMMENABLE[4], CFGINTERRUPTMSIMMENABLE_OUT[4]);
  buf B_CFGINTERRUPTMSIMMENABLE5 (CFGINTERRUPTMSIMMENABLE[5], CFGINTERRUPTMSIMMENABLE_OUT[5]);
  buf B_CFGINTERRUPTMSISENT (CFGINTERRUPTMSISENT, CFGINTERRUPTMSISENT_OUT);
  buf B_CFGINTERRUPTMSIVFENABLE0 (CFGINTERRUPTMSIVFENABLE[0], CFGINTERRUPTMSIVFENABLE_OUT[0]);
  buf B_CFGINTERRUPTMSIVFENABLE1 (CFGINTERRUPTMSIVFENABLE[1], CFGINTERRUPTMSIVFENABLE_OUT[1]);
  buf B_CFGINTERRUPTMSIVFENABLE2 (CFGINTERRUPTMSIVFENABLE[2], CFGINTERRUPTMSIVFENABLE_OUT[2]);
  buf B_CFGINTERRUPTMSIVFENABLE3 (CFGINTERRUPTMSIVFENABLE[3], CFGINTERRUPTMSIVFENABLE_OUT[3]);
  buf B_CFGINTERRUPTMSIVFENABLE4 (CFGINTERRUPTMSIVFENABLE[4], CFGINTERRUPTMSIVFENABLE_OUT[4]);
  buf B_CFGINTERRUPTMSIVFENABLE5 (CFGINTERRUPTMSIVFENABLE[5], CFGINTERRUPTMSIVFENABLE_OUT[5]);
  buf B_CFGINTERRUPTMSIXENABLE0 (CFGINTERRUPTMSIXENABLE[0], CFGINTERRUPTMSIXENABLE_OUT[0]);
  buf B_CFGINTERRUPTMSIXENABLE1 (CFGINTERRUPTMSIXENABLE[1], CFGINTERRUPTMSIXENABLE_OUT[1]);
  buf B_CFGINTERRUPTMSIXFAIL (CFGINTERRUPTMSIXFAIL, CFGINTERRUPTMSIXFAIL_OUT);
  buf B_CFGINTERRUPTMSIXMASK0 (CFGINTERRUPTMSIXMASK[0], CFGINTERRUPTMSIXMASK_OUT[0]);
  buf B_CFGINTERRUPTMSIXMASK1 (CFGINTERRUPTMSIXMASK[1], CFGINTERRUPTMSIXMASK_OUT[1]);
  buf B_CFGINTERRUPTMSIXSENT (CFGINTERRUPTMSIXSENT, CFGINTERRUPTMSIXSENT_OUT);
  buf B_CFGINTERRUPTMSIXVFENABLE0 (CFGINTERRUPTMSIXVFENABLE[0], CFGINTERRUPTMSIXVFENABLE_OUT[0]);
  buf B_CFGINTERRUPTMSIXVFENABLE1 (CFGINTERRUPTMSIXVFENABLE[1], CFGINTERRUPTMSIXVFENABLE_OUT[1]);
  buf B_CFGINTERRUPTMSIXVFENABLE2 (CFGINTERRUPTMSIXVFENABLE[2], CFGINTERRUPTMSIXVFENABLE_OUT[2]);
  buf B_CFGINTERRUPTMSIXVFENABLE3 (CFGINTERRUPTMSIXVFENABLE[3], CFGINTERRUPTMSIXVFENABLE_OUT[3]);
  buf B_CFGINTERRUPTMSIXVFENABLE4 (CFGINTERRUPTMSIXVFENABLE[4], CFGINTERRUPTMSIXVFENABLE_OUT[4]);
  buf B_CFGINTERRUPTMSIXVFENABLE5 (CFGINTERRUPTMSIXVFENABLE[5], CFGINTERRUPTMSIXVFENABLE_OUT[5]);
  buf B_CFGINTERRUPTMSIXVFMASK0 (CFGINTERRUPTMSIXVFMASK[0], CFGINTERRUPTMSIXVFMASK_OUT[0]);
  buf B_CFGINTERRUPTMSIXVFMASK1 (CFGINTERRUPTMSIXVFMASK[1], CFGINTERRUPTMSIXVFMASK_OUT[1]);
  buf B_CFGINTERRUPTMSIXVFMASK2 (CFGINTERRUPTMSIXVFMASK[2], CFGINTERRUPTMSIXVFMASK_OUT[2]);
  buf B_CFGINTERRUPTMSIXVFMASK3 (CFGINTERRUPTMSIXVFMASK[3], CFGINTERRUPTMSIXVFMASK_OUT[3]);
  buf B_CFGINTERRUPTMSIXVFMASK4 (CFGINTERRUPTMSIXVFMASK[4], CFGINTERRUPTMSIXVFMASK_OUT[4]);
  buf B_CFGINTERRUPTMSIXVFMASK5 (CFGINTERRUPTMSIXVFMASK[5], CFGINTERRUPTMSIXVFMASK_OUT[5]);
  buf B_CFGINTERRUPTSENT (CFGINTERRUPTSENT, CFGINTERRUPTSENT_OUT);
  buf B_CFGLINKPOWERSTATE0 (CFGLINKPOWERSTATE[0], CFGLINKPOWERSTATE_OUT[0]);
  buf B_CFGLINKPOWERSTATE1 (CFGLINKPOWERSTATE[1], CFGLINKPOWERSTATE_OUT[1]);
  buf B_CFGLOCALERROR (CFGLOCALERROR, CFGLOCALERROR_OUT);
  buf B_CFGLTRENABLE (CFGLTRENABLE, CFGLTRENABLE_OUT);
  buf B_CFGLTSSMSTATE0 (CFGLTSSMSTATE[0], CFGLTSSMSTATE_OUT[0]);
  buf B_CFGLTSSMSTATE1 (CFGLTSSMSTATE[1], CFGLTSSMSTATE_OUT[1]);
  buf B_CFGLTSSMSTATE2 (CFGLTSSMSTATE[2], CFGLTSSMSTATE_OUT[2]);
  buf B_CFGLTSSMSTATE3 (CFGLTSSMSTATE[3], CFGLTSSMSTATE_OUT[3]);
  buf B_CFGLTSSMSTATE4 (CFGLTSSMSTATE[4], CFGLTSSMSTATE_OUT[4]);
  buf B_CFGLTSSMSTATE5 (CFGLTSSMSTATE[5], CFGLTSSMSTATE_OUT[5]);
  buf B_CFGMAXPAYLOAD0 (CFGMAXPAYLOAD[0], CFGMAXPAYLOAD_OUT[0]);
  buf B_CFGMAXPAYLOAD1 (CFGMAXPAYLOAD[1], CFGMAXPAYLOAD_OUT[1]);
  buf B_CFGMAXPAYLOAD2 (CFGMAXPAYLOAD[2], CFGMAXPAYLOAD_OUT[2]);
  buf B_CFGMAXREADREQ0 (CFGMAXREADREQ[0], CFGMAXREADREQ_OUT[0]);
  buf B_CFGMAXREADREQ1 (CFGMAXREADREQ[1], CFGMAXREADREQ_OUT[1]);
  buf B_CFGMAXREADREQ2 (CFGMAXREADREQ[2], CFGMAXREADREQ_OUT[2]);
  buf B_CFGMCUPDATEDONE (CFGMCUPDATEDONE, CFGMCUPDATEDONE_OUT);
  buf B_CFGMGMTREADDATA0 (CFGMGMTREADDATA[0], CFGMGMTREADDATA_OUT[0]);
  buf B_CFGMGMTREADDATA1 (CFGMGMTREADDATA[1], CFGMGMTREADDATA_OUT[1]);
  buf B_CFGMGMTREADDATA10 (CFGMGMTREADDATA[10], CFGMGMTREADDATA_OUT[10]);
  buf B_CFGMGMTREADDATA11 (CFGMGMTREADDATA[11], CFGMGMTREADDATA_OUT[11]);
  buf B_CFGMGMTREADDATA12 (CFGMGMTREADDATA[12], CFGMGMTREADDATA_OUT[12]);
  buf B_CFGMGMTREADDATA13 (CFGMGMTREADDATA[13], CFGMGMTREADDATA_OUT[13]);
  buf B_CFGMGMTREADDATA14 (CFGMGMTREADDATA[14], CFGMGMTREADDATA_OUT[14]);
  buf B_CFGMGMTREADDATA15 (CFGMGMTREADDATA[15], CFGMGMTREADDATA_OUT[15]);
  buf B_CFGMGMTREADDATA16 (CFGMGMTREADDATA[16], CFGMGMTREADDATA_OUT[16]);
  buf B_CFGMGMTREADDATA17 (CFGMGMTREADDATA[17], CFGMGMTREADDATA_OUT[17]);
  buf B_CFGMGMTREADDATA18 (CFGMGMTREADDATA[18], CFGMGMTREADDATA_OUT[18]);
  buf B_CFGMGMTREADDATA19 (CFGMGMTREADDATA[19], CFGMGMTREADDATA_OUT[19]);
  buf B_CFGMGMTREADDATA2 (CFGMGMTREADDATA[2], CFGMGMTREADDATA_OUT[2]);
  buf B_CFGMGMTREADDATA20 (CFGMGMTREADDATA[20], CFGMGMTREADDATA_OUT[20]);
  buf B_CFGMGMTREADDATA21 (CFGMGMTREADDATA[21], CFGMGMTREADDATA_OUT[21]);
  buf B_CFGMGMTREADDATA22 (CFGMGMTREADDATA[22], CFGMGMTREADDATA_OUT[22]);
  buf B_CFGMGMTREADDATA23 (CFGMGMTREADDATA[23], CFGMGMTREADDATA_OUT[23]);
  buf B_CFGMGMTREADDATA24 (CFGMGMTREADDATA[24], CFGMGMTREADDATA_OUT[24]);
  buf B_CFGMGMTREADDATA25 (CFGMGMTREADDATA[25], CFGMGMTREADDATA_OUT[25]);
  buf B_CFGMGMTREADDATA26 (CFGMGMTREADDATA[26], CFGMGMTREADDATA_OUT[26]);
  buf B_CFGMGMTREADDATA27 (CFGMGMTREADDATA[27], CFGMGMTREADDATA_OUT[27]);
  buf B_CFGMGMTREADDATA28 (CFGMGMTREADDATA[28], CFGMGMTREADDATA_OUT[28]);
  buf B_CFGMGMTREADDATA29 (CFGMGMTREADDATA[29], CFGMGMTREADDATA_OUT[29]);
  buf B_CFGMGMTREADDATA3 (CFGMGMTREADDATA[3], CFGMGMTREADDATA_OUT[3]);
  buf B_CFGMGMTREADDATA30 (CFGMGMTREADDATA[30], CFGMGMTREADDATA_OUT[30]);
  buf B_CFGMGMTREADDATA31 (CFGMGMTREADDATA[31], CFGMGMTREADDATA_OUT[31]);
  buf B_CFGMGMTREADDATA4 (CFGMGMTREADDATA[4], CFGMGMTREADDATA_OUT[4]);
  buf B_CFGMGMTREADDATA5 (CFGMGMTREADDATA[5], CFGMGMTREADDATA_OUT[5]);
  buf B_CFGMGMTREADDATA6 (CFGMGMTREADDATA[6], CFGMGMTREADDATA_OUT[6]);
  buf B_CFGMGMTREADDATA7 (CFGMGMTREADDATA[7], CFGMGMTREADDATA_OUT[7]);
  buf B_CFGMGMTREADDATA8 (CFGMGMTREADDATA[8], CFGMGMTREADDATA_OUT[8]);
  buf B_CFGMGMTREADDATA9 (CFGMGMTREADDATA[9], CFGMGMTREADDATA_OUT[9]);
  buf B_CFGMGMTREADWRITEDONE (CFGMGMTREADWRITEDONE, CFGMGMTREADWRITEDONE_OUT);
  buf B_CFGMSGRECEIVED (CFGMSGRECEIVED, CFGMSGRECEIVED_OUT);
  buf B_CFGMSGRECEIVEDDATA0 (CFGMSGRECEIVEDDATA[0], CFGMSGRECEIVEDDATA_OUT[0]);
  buf B_CFGMSGRECEIVEDDATA1 (CFGMSGRECEIVEDDATA[1], CFGMSGRECEIVEDDATA_OUT[1]);
  buf B_CFGMSGRECEIVEDDATA2 (CFGMSGRECEIVEDDATA[2], CFGMSGRECEIVEDDATA_OUT[2]);
  buf B_CFGMSGRECEIVEDDATA3 (CFGMSGRECEIVEDDATA[3], CFGMSGRECEIVEDDATA_OUT[3]);
  buf B_CFGMSGRECEIVEDDATA4 (CFGMSGRECEIVEDDATA[4], CFGMSGRECEIVEDDATA_OUT[4]);
  buf B_CFGMSGRECEIVEDDATA5 (CFGMSGRECEIVEDDATA[5], CFGMSGRECEIVEDDATA_OUT[5]);
  buf B_CFGMSGRECEIVEDDATA6 (CFGMSGRECEIVEDDATA[6], CFGMSGRECEIVEDDATA_OUT[6]);
  buf B_CFGMSGRECEIVEDDATA7 (CFGMSGRECEIVEDDATA[7], CFGMSGRECEIVEDDATA_OUT[7]);
  buf B_CFGMSGRECEIVEDTYPE0 (CFGMSGRECEIVEDTYPE[0], CFGMSGRECEIVEDTYPE_OUT[0]);
  buf B_CFGMSGRECEIVEDTYPE1 (CFGMSGRECEIVEDTYPE[1], CFGMSGRECEIVEDTYPE_OUT[1]);
  buf B_CFGMSGRECEIVEDTYPE2 (CFGMSGRECEIVEDTYPE[2], CFGMSGRECEIVEDTYPE_OUT[2]);
  buf B_CFGMSGRECEIVEDTYPE3 (CFGMSGRECEIVEDTYPE[3], CFGMSGRECEIVEDTYPE_OUT[3]);
  buf B_CFGMSGRECEIVEDTYPE4 (CFGMSGRECEIVEDTYPE[4], CFGMSGRECEIVEDTYPE_OUT[4]);
  buf B_CFGMSGTRANSMITDONE (CFGMSGTRANSMITDONE, CFGMSGTRANSMITDONE_OUT);
  buf B_CFGNEGOTIATEDWIDTH0 (CFGNEGOTIATEDWIDTH[0], CFGNEGOTIATEDWIDTH_OUT[0]);
  buf B_CFGNEGOTIATEDWIDTH1 (CFGNEGOTIATEDWIDTH[1], CFGNEGOTIATEDWIDTH_OUT[1]);
  buf B_CFGNEGOTIATEDWIDTH2 (CFGNEGOTIATEDWIDTH[2], CFGNEGOTIATEDWIDTH_OUT[2]);
  buf B_CFGNEGOTIATEDWIDTH3 (CFGNEGOTIATEDWIDTH[3], CFGNEGOTIATEDWIDTH_OUT[3]);
  buf B_CFGOBFFENABLE0 (CFGOBFFENABLE[0], CFGOBFFENABLE_OUT[0]);
  buf B_CFGOBFFENABLE1 (CFGOBFFENABLE[1], CFGOBFFENABLE_OUT[1]);
  buf B_CFGPERFUNCSTATUSDATA0 (CFGPERFUNCSTATUSDATA[0], CFGPERFUNCSTATUSDATA_OUT[0]);
  buf B_CFGPERFUNCSTATUSDATA1 (CFGPERFUNCSTATUSDATA[1], CFGPERFUNCSTATUSDATA_OUT[1]);
  buf B_CFGPERFUNCSTATUSDATA10 (CFGPERFUNCSTATUSDATA[10], CFGPERFUNCSTATUSDATA_OUT[10]);
  buf B_CFGPERFUNCSTATUSDATA11 (CFGPERFUNCSTATUSDATA[11], CFGPERFUNCSTATUSDATA_OUT[11]);
  buf B_CFGPERFUNCSTATUSDATA12 (CFGPERFUNCSTATUSDATA[12], CFGPERFUNCSTATUSDATA_OUT[12]);
  buf B_CFGPERFUNCSTATUSDATA13 (CFGPERFUNCSTATUSDATA[13], CFGPERFUNCSTATUSDATA_OUT[13]);
  buf B_CFGPERFUNCSTATUSDATA14 (CFGPERFUNCSTATUSDATA[14], CFGPERFUNCSTATUSDATA_OUT[14]);
  buf B_CFGPERFUNCSTATUSDATA15 (CFGPERFUNCSTATUSDATA[15], CFGPERFUNCSTATUSDATA_OUT[15]);
  buf B_CFGPERFUNCSTATUSDATA2 (CFGPERFUNCSTATUSDATA[2], CFGPERFUNCSTATUSDATA_OUT[2]);
  buf B_CFGPERFUNCSTATUSDATA3 (CFGPERFUNCSTATUSDATA[3], CFGPERFUNCSTATUSDATA_OUT[3]);
  buf B_CFGPERFUNCSTATUSDATA4 (CFGPERFUNCSTATUSDATA[4], CFGPERFUNCSTATUSDATA_OUT[4]);
  buf B_CFGPERFUNCSTATUSDATA5 (CFGPERFUNCSTATUSDATA[5], CFGPERFUNCSTATUSDATA_OUT[5]);
  buf B_CFGPERFUNCSTATUSDATA6 (CFGPERFUNCSTATUSDATA[6], CFGPERFUNCSTATUSDATA_OUT[6]);
  buf B_CFGPERFUNCSTATUSDATA7 (CFGPERFUNCSTATUSDATA[7], CFGPERFUNCSTATUSDATA_OUT[7]);
  buf B_CFGPERFUNCSTATUSDATA8 (CFGPERFUNCSTATUSDATA[8], CFGPERFUNCSTATUSDATA_OUT[8]);
  buf B_CFGPERFUNCSTATUSDATA9 (CFGPERFUNCSTATUSDATA[9], CFGPERFUNCSTATUSDATA_OUT[9]);
  buf B_CFGPERFUNCTIONUPDATEDONE (CFGPERFUNCTIONUPDATEDONE, CFGPERFUNCTIONUPDATEDONE_OUT);
  buf B_CFGPHYLINKDOWN (CFGPHYLINKDOWN, CFGPHYLINKDOWN_OUT);
  buf B_CFGPHYLINKSTATUS0 (CFGPHYLINKSTATUS[0], CFGPHYLINKSTATUS_OUT[0]);
  buf B_CFGPHYLINKSTATUS1 (CFGPHYLINKSTATUS[1], CFGPHYLINKSTATUS_OUT[1]);
  buf B_CFGPLSTATUSCHANGE (CFGPLSTATUSCHANGE, CFGPLSTATUSCHANGE_OUT);
  buf B_CFGPOWERSTATECHANGEINTERRUPT (CFGPOWERSTATECHANGEINTERRUPT, CFGPOWERSTATECHANGEINTERRUPT_OUT);
  buf B_CFGRCBSTATUS0 (CFGRCBSTATUS[0], CFGRCBSTATUS_OUT[0]);
  buf B_CFGRCBSTATUS1 (CFGRCBSTATUS[1], CFGRCBSTATUS_OUT[1]);
  buf B_CFGTPHFUNCTIONNUM0 (CFGTPHFUNCTIONNUM[0], CFGTPHFUNCTIONNUM_OUT[0]);
  buf B_CFGTPHFUNCTIONNUM1 (CFGTPHFUNCTIONNUM[1], CFGTPHFUNCTIONNUM_OUT[1]);
  buf B_CFGTPHFUNCTIONNUM2 (CFGTPHFUNCTIONNUM[2], CFGTPHFUNCTIONNUM_OUT[2]);
  buf B_CFGTPHREQUESTERENABLE0 (CFGTPHREQUESTERENABLE[0], CFGTPHREQUESTERENABLE_OUT[0]);
  buf B_CFGTPHREQUESTERENABLE1 (CFGTPHREQUESTERENABLE[1], CFGTPHREQUESTERENABLE_OUT[1]);
  buf B_CFGTPHSTMODE0 (CFGTPHSTMODE[0], CFGTPHSTMODE_OUT[0]);
  buf B_CFGTPHSTMODE1 (CFGTPHSTMODE[1], CFGTPHSTMODE_OUT[1]);
  buf B_CFGTPHSTMODE2 (CFGTPHSTMODE[2], CFGTPHSTMODE_OUT[2]);
  buf B_CFGTPHSTMODE3 (CFGTPHSTMODE[3], CFGTPHSTMODE_OUT[3]);
  buf B_CFGTPHSTMODE4 (CFGTPHSTMODE[4], CFGTPHSTMODE_OUT[4]);
  buf B_CFGTPHSTMODE5 (CFGTPHSTMODE[5], CFGTPHSTMODE_OUT[5]);
  buf B_CFGTPHSTTADDRESS0 (CFGTPHSTTADDRESS[0], CFGTPHSTTADDRESS_OUT[0]);
  buf B_CFGTPHSTTADDRESS1 (CFGTPHSTTADDRESS[1], CFGTPHSTTADDRESS_OUT[1]);
  buf B_CFGTPHSTTADDRESS2 (CFGTPHSTTADDRESS[2], CFGTPHSTTADDRESS_OUT[2]);
  buf B_CFGTPHSTTADDRESS3 (CFGTPHSTTADDRESS[3], CFGTPHSTTADDRESS_OUT[3]);
  buf B_CFGTPHSTTADDRESS4 (CFGTPHSTTADDRESS[4], CFGTPHSTTADDRESS_OUT[4]);
  buf B_CFGTPHSTTREADENABLE (CFGTPHSTTREADENABLE, CFGTPHSTTREADENABLE_OUT);
  buf B_CFGTPHSTTWRITEBYTEVALID0 (CFGTPHSTTWRITEBYTEVALID[0], CFGTPHSTTWRITEBYTEVALID_OUT[0]);
  buf B_CFGTPHSTTWRITEBYTEVALID1 (CFGTPHSTTWRITEBYTEVALID[1], CFGTPHSTTWRITEBYTEVALID_OUT[1]);
  buf B_CFGTPHSTTWRITEBYTEVALID2 (CFGTPHSTTWRITEBYTEVALID[2], CFGTPHSTTWRITEBYTEVALID_OUT[2]);
  buf B_CFGTPHSTTWRITEBYTEVALID3 (CFGTPHSTTWRITEBYTEVALID[3], CFGTPHSTTWRITEBYTEVALID_OUT[3]);
  buf B_CFGTPHSTTWRITEDATA0 (CFGTPHSTTWRITEDATA[0], CFGTPHSTTWRITEDATA_OUT[0]);
  buf B_CFGTPHSTTWRITEDATA1 (CFGTPHSTTWRITEDATA[1], CFGTPHSTTWRITEDATA_OUT[1]);
  buf B_CFGTPHSTTWRITEDATA10 (CFGTPHSTTWRITEDATA[10], CFGTPHSTTWRITEDATA_OUT[10]);
  buf B_CFGTPHSTTWRITEDATA11 (CFGTPHSTTWRITEDATA[11], CFGTPHSTTWRITEDATA_OUT[11]);
  buf B_CFGTPHSTTWRITEDATA12 (CFGTPHSTTWRITEDATA[12], CFGTPHSTTWRITEDATA_OUT[12]);
  buf B_CFGTPHSTTWRITEDATA13 (CFGTPHSTTWRITEDATA[13], CFGTPHSTTWRITEDATA_OUT[13]);
  buf B_CFGTPHSTTWRITEDATA14 (CFGTPHSTTWRITEDATA[14], CFGTPHSTTWRITEDATA_OUT[14]);
  buf B_CFGTPHSTTWRITEDATA15 (CFGTPHSTTWRITEDATA[15], CFGTPHSTTWRITEDATA_OUT[15]);
  buf B_CFGTPHSTTWRITEDATA16 (CFGTPHSTTWRITEDATA[16], CFGTPHSTTWRITEDATA_OUT[16]);
  buf B_CFGTPHSTTWRITEDATA17 (CFGTPHSTTWRITEDATA[17], CFGTPHSTTWRITEDATA_OUT[17]);
  buf B_CFGTPHSTTWRITEDATA18 (CFGTPHSTTWRITEDATA[18], CFGTPHSTTWRITEDATA_OUT[18]);
  buf B_CFGTPHSTTWRITEDATA19 (CFGTPHSTTWRITEDATA[19], CFGTPHSTTWRITEDATA_OUT[19]);
  buf B_CFGTPHSTTWRITEDATA2 (CFGTPHSTTWRITEDATA[2], CFGTPHSTTWRITEDATA_OUT[2]);
  buf B_CFGTPHSTTWRITEDATA20 (CFGTPHSTTWRITEDATA[20], CFGTPHSTTWRITEDATA_OUT[20]);
  buf B_CFGTPHSTTWRITEDATA21 (CFGTPHSTTWRITEDATA[21], CFGTPHSTTWRITEDATA_OUT[21]);
  buf B_CFGTPHSTTWRITEDATA22 (CFGTPHSTTWRITEDATA[22], CFGTPHSTTWRITEDATA_OUT[22]);
  buf B_CFGTPHSTTWRITEDATA23 (CFGTPHSTTWRITEDATA[23], CFGTPHSTTWRITEDATA_OUT[23]);
  buf B_CFGTPHSTTWRITEDATA24 (CFGTPHSTTWRITEDATA[24], CFGTPHSTTWRITEDATA_OUT[24]);
  buf B_CFGTPHSTTWRITEDATA25 (CFGTPHSTTWRITEDATA[25], CFGTPHSTTWRITEDATA_OUT[25]);
  buf B_CFGTPHSTTWRITEDATA26 (CFGTPHSTTWRITEDATA[26], CFGTPHSTTWRITEDATA_OUT[26]);
  buf B_CFGTPHSTTWRITEDATA27 (CFGTPHSTTWRITEDATA[27], CFGTPHSTTWRITEDATA_OUT[27]);
  buf B_CFGTPHSTTWRITEDATA28 (CFGTPHSTTWRITEDATA[28], CFGTPHSTTWRITEDATA_OUT[28]);
  buf B_CFGTPHSTTWRITEDATA29 (CFGTPHSTTWRITEDATA[29], CFGTPHSTTWRITEDATA_OUT[29]);
  buf B_CFGTPHSTTWRITEDATA3 (CFGTPHSTTWRITEDATA[3], CFGTPHSTTWRITEDATA_OUT[3]);
  buf B_CFGTPHSTTWRITEDATA30 (CFGTPHSTTWRITEDATA[30], CFGTPHSTTWRITEDATA_OUT[30]);
  buf B_CFGTPHSTTWRITEDATA31 (CFGTPHSTTWRITEDATA[31], CFGTPHSTTWRITEDATA_OUT[31]);
  buf B_CFGTPHSTTWRITEDATA4 (CFGTPHSTTWRITEDATA[4], CFGTPHSTTWRITEDATA_OUT[4]);
  buf B_CFGTPHSTTWRITEDATA5 (CFGTPHSTTWRITEDATA[5], CFGTPHSTTWRITEDATA_OUT[5]);
  buf B_CFGTPHSTTWRITEDATA6 (CFGTPHSTTWRITEDATA[6], CFGTPHSTTWRITEDATA_OUT[6]);
  buf B_CFGTPHSTTWRITEDATA7 (CFGTPHSTTWRITEDATA[7], CFGTPHSTTWRITEDATA_OUT[7]);
  buf B_CFGTPHSTTWRITEDATA8 (CFGTPHSTTWRITEDATA[8], CFGTPHSTTWRITEDATA_OUT[8]);
  buf B_CFGTPHSTTWRITEDATA9 (CFGTPHSTTWRITEDATA[9], CFGTPHSTTWRITEDATA_OUT[9]);
  buf B_CFGTPHSTTWRITEENABLE (CFGTPHSTTWRITEENABLE, CFGTPHSTTWRITEENABLE_OUT);
  buf B_CFGVFFLRINPROCESS0 (CFGVFFLRINPROCESS[0], CFGVFFLRINPROCESS_OUT[0]);
  buf B_CFGVFFLRINPROCESS1 (CFGVFFLRINPROCESS[1], CFGVFFLRINPROCESS_OUT[1]);
  buf B_CFGVFFLRINPROCESS2 (CFGVFFLRINPROCESS[2], CFGVFFLRINPROCESS_OUT[2]);
  buf B_CFGVFFLRINPROCESS3 (CFGVFFLRINPROCESS[3], CFGVFFLRINPROCESS_OUT[3]);
  buf B_CFGVFFLRINPROCESS4 (CFGVFFLRINPROCESS[4], CFGVFFLRINPROCESS_OUT[4]);
  buf B_CFGVFFLRINPROCESS5 (CFGVFFLRINPROCESS[5], CFGVFFLRINPROCESS_OUT[5]);
  buf B_CFGVFPOWERSTATE0 (CFGVFPOWERSTATE[0], CFGVFPOWERSTATE_OUT[0]);
  buf B_CFGVFPOWERSTATE1 (CFGVFPOWERSTATE[1], CFGVFPOWERSTATE_OUT[1]);
  buf B_CFGVFPOWERSTATE10 (CFGVFPOWERSTATE[10], CFGVFPOWERSTATE_OUT[10]);
  buf B_CFGVFPOWERSTATE11 (CFGVFPOWERSTATE[11], CFGVFPOWERSTATE_OUT[11]);
  buf B_CFGVFPOWERSTATE12 (CFGVFPOWERSTATE[12], CFGVFPOWERSTATE_OUT[12]);
  buf B_CFGVFPOWERSTATE13 (CFGVFPOWERSTATE[13], CFGVFPOWERSTATE_OUT[13]);
  buf B_CFGVFPOWERSTATE14 (CFGVFPOWERSTATE[14], CFGVFPOWERSTATE_OUT[14]);
  buf B_CFGVFPOWERSTATE15 (CFGVFPOWERSTATE[15], CFGVFPOWERSTATE_OUT[15]);
  buf B_CFGVFPOWERSTATE16 (CFGVFPOWERSTATE[16], CFGVFPOWERSTATE_OUT[16]);
  buf B_CFGVFPOWERSTATE17 (CFGVFPOWERSTATE[17], CFGVFPOWERSTATE_OUT[17]);
  buf B_CFGVFPOWERSTATE2 (CFGVFPOWERSTATE[2], CFGVFPOWERSTATE_OUT[2]);
  buf B_CFGVFPOWERSTATE3 (CFGVFPOWERSTATE[3], CFGVFPOWERSTATE_OUT[3]);
  buf B_CFGVFPOWERSTATE4 (CFGVFPOWERSTATE[4], CFGVFPOWERSTATE_OUT[4]);
  buf B_CFGVFPOWERSTATE5 (CFGVFPOWERSTATE[5], CFGVFPOWERSTATE_OUT[5]);
  buf B_CFGVFPOWERSTATE6 (CFGVFPOWERSTATE[6], CFGVFPOWERSTATE_OUT[6]);
  buf B_CFGVFPOWERSTATE7 (CFGVFPOWERSTATE[7], CFGVFPOWERSTATE_OUT[7]);
  buf B_CFGVFPOWERSTATE8 (CFGVFPOWERSTATE[8], CFGVFPOWERSTATE_OUT[8]);
  buf B_CFGVFPOWERSTATE9 (CFGVFPOWERSTATE[9], CFGVFPOWERSTATE_OUT[9]);
  buf B_CFGVFSTATUS0 (CFGVFSTATUS[0], CFGVFSTATUS_OUT[0]);
  buf B_CFGVFSTATUS1 (CFGVFSTATUS[1], CFGVFSTATUS_OUT[1]);
  buf B_CFGVFSTATUS10 (CFGVFSTATUS[10], CFGVFSTATUS_OUT[10]);
  buf B_CFGVFSTATUS11 (CFGVFSTATUS[11], CFGVFSTATUS_OUT[11]);
  buf B_CFGVFSTATUS2 (CFGVFSTATUS[2], CFGVFSTATUS_OUT[2]);
  buf B_CFGVFSTATUS3 (CFGVFSTATUS[3], CFGVFSTATUS_OUT[3]);
  buf B_CFGVFSTATUS4 (CFGVFSTATUS[4], CFGVFSTATUS_OUT[4]);
  buf B_CFGVFSTATUS5 (CFGVFSTATUS[5], CFGVFSTATUS_OUT[5]);
  buf B_CFGVFSTATUS6 (CFGVFSTATUS[6], CFGVFSTATUS_OUT[6]);
  buf B_CFGVFSTATUS7 (CFGVFSTATUS[7], CFGVFSTATUS_OUT[7]);
  buf B_CFGVFSTATUS8 (CFGVFSTATUS[8], CFGVFSTATUS_OUT[8]);
  buf B_CFGVFSTATUS9 (CFGVFSTATUS[9], CFGVFSTATUS_OUT[9]);
  buf B_CFGVFTPHREQUESTERENABLE0 (CFGVFTPHREQUESTERENABLE[0], CFGVFTPHREQUESTERENABLE_OUT[0]);
  buf B_CFGVFTPHREQUESTERENABLE1 (CFGVFTPHREQUESTERENABLE[1], CFGVFTPHREQUESTERENABLE_OUT[1]);
  buf B_CFGVFTPHREQUESTERENABLE2 (CFGVFTPHREQUESTERENABLE[2], CFGVFTPHREQUESTERENABLE_OUT[2]);
  buf B_CFGVFTPHREQUESTERENABLE3 (CFGVFTPHREQUESTERENABLE[3], CFGVFTPHREQUESTERENABLE_OUT[3]);
  buf B_CFGVFTPHREQUESTERENABLE4 (CFGVFTPHREQUESTERENABLE[4], CFGVFTPHREQUESTERENABLE_OUT[4]);
  buf B_CFGVFTPHREQUESTERENABLE5 (CFGVFTPHREQUESTERENABLE[5], CFGVFTPHREQUESTERENABLE_OUT[5]);
  buf B_CFGVFTPHSTMODE0 (CFGVFTPHSTMODE[0], CFGVFTPHSTMODE_OUT[0]);
  buf B_CFGVFTPHSTMODE1 (CFGVFTPHSTMODE[1], CFGVFTPHSTMODE_OUT[1]);
  buf B_CFGVFTPHSTMODE10 (CFGVFTPHSTMODE[10], CFGVFTPHSTMODE_OUT[10]);
  buf B_CFGVFTPHSTMODE11 (CFGVFTPHSTMODE[11], CFGVFTPHSTMODE_OUT[11]);
  buf B_CFGVFTPHSTMODE12 (CFGVFTPHSTMODE[12], CFGVFTPHSTMODE_OUT[12]);
  buf B_CFGVFTPHSTMODE13 (CFGVFTPHSTMODE[13], CFGVFTPHSTMODE_OUT[13]);
  buf B_CFGVFTPHSTMODE14 (CFGVFTPHSTMODE[14], CFGVFTPHSTMODE_OUT[14]);
  buf B_CFGVFTPHSTMODE15 (CFGVFTPHSTMODE[15], CFGVFTPHSTMODE_OUT[15]);
  buf B_CFGVFTPHSTMODE16 (CFGVFTPHSTMODE[16], CFGVFTPHSTMODE_OUT[16]);
  buf B_CFGVFTPHSTMODE17 (CFGVFTPHSTMODE[17], CFGVFTPHSTMODE_OUT[17]);
  buf B_CFGVFTPHSTMODE2 (CFGVFTPHSTMODE[2], CFGVFTPHSTMODE_OUT[2]);
  buf B_CFGVFTPHSTMODE3 (CFGVFTPHSTMODE[3], CFGVFTPHSTMODE_OUT[3]);
  buf B_CFGVFTPHSTMODE4 (CFGVFTPHSTMODE[4], CFGVFTPHSTMODE_OUT[4]);
  buf B_CFGVFTPHSTMODE5 (CFGVFTPHSTMODE[5], CFGVFTPHSTMODE_OUT[5]);
  buf B_CFGVFTPHSTMODE6 (CFGVFTPHSTMODE[6], CFGVFTPHSTMODE_OUT[6]);
  buf B_CFGVFTPHSTMODE7 (CFGVFTPHSTMODE[7], CFGVFTPHSTMODE_OUT[7]);
  buf B_CFGVFTPHSTMODE8 (CFGVFTPHSTMODE[8], CFGVFTPHSTMODE_OUT[8]);
  buf B_CFGVFTPHSTMODE9 (CFGVFTPHSTMODE[9], CFGVFTPHSTMODE_OUT[9]);
  buf B_DBGDATAOUT0 (DBGDATAOUT[0], DBGDATAOUT_OUT[0]);
  buf B_DBGDATAOUT1 (DBGDATAOUT[1], DBGDATAOUT_OUT[1]);
  buf B_DBGDATAOUT10 (DBGDATAOUT[10], DBGDATAOUT_OUT[10]);
  buf B_DBGDATAOUT11 (DBGDATAOUT[11], DBGDATAOUT_OUT[11]);
  buf B_DBGDATAOUT12 (DBGDATAOUT[12], DBGDATAOUT_OUT[12]);
  buf B_DBGDATAOUT13 (DBGDATAOUT[13], DBGDATAOUT_OUT[13]);
  buf B_DBGDATAOUT14 (DBGDATAOUT[14], DBGDATAOUT_OUT[14]);
  buf B_DBGDATAOUT15 (DBGDATAOUT[15], DBGDATAOUT_OUT[15]);
  buf B_DBGDATAOUT2 (DBGDATAOUT[2], DBGDATAOUT_OUT[2]);
  buf B_DBGDATAOUT3 (DBGDATAOUT[3], DBGDATAOUT_OUT[3]);
  buf B_DBGDATAOUT4 (DBGDATAOUT[4], DBGDATAOUT_OUT[4]);
  buf B_DBGDATAOUT5 (DBGDATAOUT[5], DBGDATAOUT_OUT[5]);
  buf B_DBGDATAOUT6 (DBGDATAOUT[6], DBGDATAOUT_OUT[6]);
  buf B_DBGDATAOUT7 (DBGDATAOUT[7], DBGDATAOUT_OUT[7]);
  buf B_DBGDATAOUT8 (DBGDATAOUT[8], DBGDATAOUT_OUT[8]);
  buf B_DBGDATAOUT9 (DBGDATAOUT[9], DBGDATAOUT_OUT[9]);
  buf B_DRPDO0 (DRPDO[0], DRPDO_OUT[0]);
  buf B_DRPDO1 (DRPDO[1], DRPDO_OUT[1]);
  buf B_DRPDO10 (DRPDO[10], DRPDO_OUT[10]);
  buf B_DRPDO11 (DRPDO[11], DRPDO_OUT[11]);
  buf B_DRPDO12 (DRPDO[12], DRPDO_OUT[12]);
  buf B_DRPDO13 (DRPDO[13], DRPDO_OUT[13]);
  buf B_DRPDO14 (DRPDO[14], DRPDO_OUT[14]);
  buf B_DRPDO15 (DRPDO[15], DRPDO_OUT[15]);
  buf B_DRPDO2 (DRPDO[2], DRPDO_OUT[2]);
  buf B_DRPDO3 (DRPDO[3], DRPDO_OUT[3]);
  buf B_DRPDO4 (DRPDO[4], DRPDO_OUT[4]);
  buf B_DRPDO5 (DRPDO[5], DRPDO_OUT[5]);
  buf B_DRPDO6 (DRPDO[6], DRPDO_OUT[6]);
  buf B_DRPDO7 (DRPDO[7], DRPDO_OUT[7]);
  buf B_DRPDO8 (DRPDO[8], DRPDO_OUT[8]);
  buf B_DRPDO9 (DRPDO[9], DRPDO_OUT[9]);
  buf B_DRPRDY (DRPRDY, DRPRDY_OUT);
  buf B_MAXISCQTDATA0 (MAXISCQTDATA[0], MAXISCQTDATA_OUT[0]);
  buf B_MAXISCQTDATA1 (MAXISCQTDATA[1], MAXISCQTDATA_OUT[1]);
  buf B_MAXISCQTDATA10 (MAXISCQTDATA[10], MAXISCQTDATA_OUT[10]);
  buf B_MAXISCQTDATA100 (MAXISCQTDATA[100], MAXISCQTDATA_OUT[100]);
  buf B_MAXISCQTDATA101 (MAXISCQTDATA[101], MAXISCQTDATA_OUT[101]);
  buf B_MAXISCQTDATA102 (MAXISCQTDATA[102], MAXISCQTDATA_OUT[102]);
  buf B_MAXISCQTDATA103 (MAXISCQTDATA[103], MAXISCQTDATA_OUT[103]);
  buf B_MAXISCQTDATA104 (MAXISCQTDATA[104], MAXISCQTDATA_OUT[104]);
  buf B_MAXISCQTDATA105 (MAXISCQTDATA[105], MAXISCQTDATA_OUT[105]);
  buf B_MAXISCQTDATA106 (MAXISCQTDATA[106], MAXISCQTDATA_OUT[106]);
  buf B_MAXISCQTDATA107 (MAXISCQTDATA[107], MAXISCQTDATA_OUT[107]);
  buf B_MAXISCQTDATA108 (MAXISCQTDATA[108], MAXISCQTDATA_OUT[108]);
  buf B_MAXISCQTDATA109 (MAXISCQTDATA[109], MAXISCQTDATA_OUT[109]);
  buf B_MAXISCQTDATA11 (MAXISCQTDATA[11], MAXISCQTDATA_OUT[11]);
  buf B_MAXISCQTDATA110 (MAXISCQTDATA[110], MAXISCQTDATA_OUT[110]);
  buf B_MAXISCQTDATA111 (MAXISCQTDATA[111], MAXISCQTDATA_OUT[111]);
  buf B_MAXISCQTDATA112 (MAXISCQTDATA[112], MAXISCQTDATA_OUT[112]);
  buf B_MAXISCQTDATA113 (MAXISCQTDATA[113], MAXISCQTDATA_OUT[113]);
  buf B_MAXISCQTDATA114 (MAXISCQTDATA[114], MAXISCQTDATA_OUT[114]);
  buf B_MAXISCQTDATA115 (MAXISCQTDATA[115], MAXISCQTDATA_OUT[115]);
  buf B_MAXISCQTDATA116 (MAXISCQTDATA[116], MAXISCQTDATA_OUT[116]);
  buf B_MAXISCQTDATA117 (MAXISCQTDATA[117], MAXISCQTDATA_OUT[117]);
  buf B_MAXISCQTDATA118 (MAXISCQTDATA[118], MAXISCQTDATA_OUT[118]);
  buf B_MAXISCQTDATA119 (MAXISCQTDATA[119], MAXISCQTDATA_OUT[119]);
  buf B_MAXISCQTDATA12 (MAXISCQTDATA[12], MAXISCQTDATA_OUT[12]);
  buf B_MAXISCQTDATA120 (MAXISCQTDATA[120], MAXISCQTDATA_OUT[120]);
  buf B_MAXISCQTDATA121 (MAXISCQTDATA[121], MAXISCQTDATA_OUT[121]);
  buf B_MAXISCQTDATA122 (MAXISCQTDATA[122], MAXISCQTDATA_OUT[122]);
  buf B_MAXISCQTDATA123 (MAXISCQTDATA[123], MAXISCQTDATA_OUT[123]);
  buf B_MAXISCQTDATA124 (MAXISCQTDATA[124], MAXISCQTDATA_OUT[124]);
  buf B_MAXISCQTDATA125 (MAXISCQTDATA[125], MAXISCQTDATA_OUT[125]);
  buf B_MAXISCQTDATA126 (MAXISCQTDATA[126], MAXISCQTDATA_OUT[126]);
  buf B_MAXISCQTDATA127 (MAXISCQTDATA[127], MAXISCQTDATA_OUT[127]);
  buf B_MAXISCQTDATA128 (MAXISCQTDATA[128], MAXISCQTDATA_OUT[128]);
  buf B_MAXISCQTDATA129 (MAXISCQTDATA[129], MAXISCQTDATA_OUT[129]);
  buf B_MAXISCQTDATA13 (MAXISCQTDATA[13], MAXISCQTDATA_OUT[13]);
  buf B_MAXISCQTDATA130 (MAXISCQTDATA[130], MAXISCQTDATA_OUT[130]);
  buf B_MAXISCQTDATA131 (MAXISCQTDATA[131], MAXISCQTDATA_OUT[131]);
  buf B_MAXISCQTDATA132 (MAXISCQTDATA[132], MAXISCQTDATA_OUT[132]);
  buf B_MAXISCQTDATA133 (MAXISCQTDATA[133], MAXISCQTDATA_OUT[133]);
  buf B_MAXISCQTDATA134 (MAXISCQTDATA[134], MAXISCQTDATA_OUT[134]);
  buf B_MAXISCQTDATA135 (MAXISCQTDATA[135], MAXISCQTDATA_OUT[135]);
  buf B_MAXISCQTDATA136 (MAXISCQTDATA[136], MAXISCQTDATA_OUT[136]);
  buf B_MAXISCQTDATA137 (MAXISCQTDATA[137], MAXISCQTDATA_OUT[137]);
  buf B_MAXISCQTDATA138 (MAXISCQTDATA[138], MAXISCQTDATA_OUT[138]);
  buf B_MAXISCQTDATA139 (MAXISCQTDATA[139], MAXISCQTDATA_OUT[139]);
  buf B_MAXISCQTDATA14 (MAXISCQTDATA[14], MAXISCQTDATA_OUT[14]);
  buf B_MAXISCQTDATA140 (MAXISCQTDATA[140], MAXISCQTDATA_OUT[140]);
  buf B_MAXISCQTDATA141 (MAXISCQTDATA[141], MAXISCQTDATA_OUT[141]);
  buf B_MAXISCQTDATA142 (MAXISCQTDATA[142], MAXISCQTDATA_OUT[142]);
  buf B_MAXISCQTDATA143 (MAXISCQTDATA[143], MAXISCQTDATA_OUT[143]);
  buf B_MAXISCQTDATA144 (MAXISCQTDATA[144], MAXISCQTDATA_OUT[144]);
  buf B_MAXISCQTDATA145 (MAXISCQTDATA[145], MAXISCQTDATA_OUT[145]);
  buf B_MAXISCQTDATA146 (MAXISCQTDATA[146], MAXISCQTDATA_OUT[146]);
  buf B_MAXISCQTDATA147 (MAXISCQTDATA[147], MAXISCQTDATA_OUT[147]);
  buf B_MAXISCQTDATA148 (MAXISCQTDATA[148], MAXISCQTDATA_OUT[148]);
  buf B_MAXISCQTDATA149 (MAXISCQTDATA[149], MAXISCQTDATA_OUT[149]);
  buf B_MAXISCQTDATA15 (MAXISCQTDATA[15], MAXISCQTDATA_OUT[15]);
  buf B_MAXISCQTDATA150 (MAXISCQTDATA[150], MAXISCQTDATA_OUT[150]);
  buf B_MAXISCQTDATA151 (MAXISCQTDATA[151], MAXISCQTDATA_OUT[151]);
  buf B_MAXISCQTDATA152 (MAXISCQTDATA[152], MAXISCQTDATA_OUT[152]);
  buf B_MAXISCQTDATA153 (MAXISCQTDATA[153], MAXISCQTDATA_OUT[153]);
  buf B_MAXISCQTDATA154 (MAXISCQTDATA[154], MAXISCQTDATA_OUT[154]);
  buf B_MAXISCQTDATA155 (MAXISCQTDATA[155], MAXISCQTDATA_OUT[155]);
  buf B_MAXISCQTDATA156 (MAXISCQTDATA[156], MAXISCQTDATA_OUT[156]);
  buf B_MAXISCQTDATA157 (MAXISCQTDATA[157], MAXISCQTDATA_OUT[157]);
  buf B_MAXISCQTDATA158 (MAXISCQTDATA[158], MAXISCQTDATA_OUT[158]);
  buf B_MAXISCQTDATA159 (MAXISCQTDATA[159], MAXISCQTDATA_OUT[159]);
  buf B_MAXISCQTDATA16 (MAXISCQTDATA[16], MAXISCQTDATA_OUT[16]);
  buf B_MAXISCQTDATA160 (MAXISCQTDATA[160], MAXISCQTDATA_OUT[160]);
  buf B_MAXISCQTDATA161 (MAXISCQTDATA[161], MAXISCQTDATA_OUT[161]);
  buf B_MAXISCQTDATA162 (MAXISCQTDATA[162], MAXISCQTDATA_OUT[162]);
  buf B_MAXISCQTDATA163 (MAXISCQTDATA[163], MAXISCQTDATA_OUT[163]);
  buf B_MAXISCQTDATA164 (MAXISCQTDATA[164], MAXISCQTDATA_OUT[164]);
  buf B_MAXISCQTDATA165 (MAXISCQTDATA[165], MAXISCQTDATA_OUT[165]);
  buf B_MAXISCQTDATA166 (MAXISCQTDATA[166], MAXISCQTDATA_OUT[166]);
  buf B_MAXISCQTDATA167 (MAXISCQTDATA[167], MAXISCQTDATA_OUT[167]);
  buf B_MAXISCQTDATA168 (MAXISCQTDATA[168], MAXISCQTDATA_OUT[168]);
  buf B_MAXISCQTDATA169 (MAXISCQTDATA[169], MAXISCQTDATA_OUT[169]);
  buf B_MAXISCQTDATA17 (MAXISCQTDATA[17], MAXISCQTDATA_OUT[17]);
  buf B_MAXISCQTDATA170 (MAXISCQTDATA[170], MAXISCQTDATA_OUT[170]);
  buf B_MAXISCQTDATA171 (MAXISCQTDATA[171], MAXISCQTDATA_OUT[171]);
  buf B_MAXISCQTDATA172 (MAXISCQTDATA[172], MAXISCQTDATA_OUT[172]);
  buf B_MAXISCQTDATA173 (MAXISCQTDATA[173], MAXISCQTDATA_OUT[173]);
  buf B_MAXISCQTDATA174 (MAXISCQTDATA[174], MAXISCQTDATA_OUT[174]);
  buf B_MAXISCQTDATA175 (MAXISCQTDATA[175], MAXISCQTDATA_OUT[175]);
  buf B_MAXISCQTDATA176 (MAXISCQTDATA[176], MAXISCQTDATA_OUT[176]);
  buf B_MAXISCQTDATA177 (MAXISCQTDATA[177], MAXISCQTDATA_OUT[177]);
  buf B_MAXISCQTDATA178 (MAXISCQTDATA[178], MAXISCQTDATA_OUT[178]);
  buf B_MAXISCQTDATA179 (MAXISCQTDATA[179], MAXISCQTDATA_OUT[179]);
  buf B_MAXISCQTDATA18 (MAXISCQTDATA[18], MAXISCQTDATA_OUT[18]);
  buf B_MAXISCQTDATA180 (MAXISCQTDATA[180], MAXISCQTDATA_OUT[180]);
  buf B_MAXISCQTDATA181 (MAXISCQTDATA[181], MAXISCQTDATA_OUT[181]);
  buf B_MAXISCQTDATA182 (MAXISCQTDATA[182], MAXISCQTDATA_OUT[182]);
  buf B_MAXISCQTDATA183 (MAXISCQTDATA[183], MAXISCQTDATA_OUT[183]);
  buf B_MAXISCQTDATA184 (MAXISCQTDATA[184], MAXISCQTDATA_OUT[184]);
  buf B_MAXISCQTDATA185 (MAXISCQTDATA[185], MAXISCQTDATA_OUT[185]);
  buf B_MAXISCQTDATA186 (MAXISCQTDATA[186], MAXISCQTDATA_OUT[186]);
  buf B_MAXISCQTDATA187 (MAXISCQTDATA[187], MAXISCQTDATA_OUT[187]);
  buf B_MAXISCQTDATA188 (MAXISCQTDATA[188], MAXISCQTDATA_OUT[188]);
  buf B_MAXISCQTDATA189 (MAXISCQTDATA[189], MAXISCQTDATA_OUT[189]);
  buf B_MAXISCQTDATA19 (MAXISCQTDATA[19], MAXISCQTDATA_OUT[19]);
  buf B_MAXISCQTDATA190 (MAXISCQTDATA[190], MAXISCQTDATA_OUT[190]);
  buf B_MAXISCQTDATA191 (MAXISCQTDATA[191], MAXISCQTDATA_OUT[191]);
  buf B_MAXISCQTDATA192 (MAXISCQTDATA[192], MAXISCQTDATA_OUT[192]);
  buf B_MAXISCQTDATA193 (MAXISCQTDATA[193], MAXISCQTDATA_OUT[193]);
  buf B_MAXISCQTDATA194 (MAXISCQTDATA[194], MAXISCQTDATA_OUT[194]);
  buf B_MAXISCQTDATA195 (MAXISCQTDATA[195], MAXISCQTDATA_OUT[195]);
  buf B_MAXISCQTDATA196 (MAXISCQTDATA[196], MAXISCQTDATA_OUT[196]);
  buf B_MAXISCQTDATA197 (MAXISCQTDATA[197], MAXISCQTDATA_OUT[197]);
  buf B_MAXISCQTDATA198 (MAXISCQTDATA[198], MAXISCQTDATA_OUT[198]);
  buf B_MAXISCQTDATA199 (MAXISCQTDATA[199], MAXISCQTDATA_OUT[199]);
  buf B_MAXISCQTDATA2 (MAXISCQTDATA[2], MAXISCQTDATA_OUT[2]);
  buf B_MAXISCQTDATA20 (MAXISCQTDATA[20], MAXISCQTDATA_OUT[20]);
  buf B_MAXISCQTDATA200 (MAXISCQTDATA[200], MAXISCQTDATA_OUT[200]);
  buf B_MAXISCQTDATA201 (MAXISCQTDATA[201], MAXISCQTDATA_OUT[201]);
  buf B_MAXISCQTDATA202 (MAXISCQTDATA[202], MAXISCQTDATA_OUT[202]);
  buf B_MAXISCQTDATA203 (MAXISCQTDATA[203], MAXISCQTDATA_OUT[203]);
  buf B_MAXISCQTDATA204 (MAXISCQTDATA[204], MAXISCQTDATA_OUT[204]);
  buf B_MAXISCQTDATA205 (MAXISCQTDATA[205], MAXISCQTDATA_OUT[205]);
  buf B_MAXISCQTDATA206 (MAXISCQTDATA[206], MAXISCQTDATA_OUT[206]);
  buf B_MAXISCQTDATA207 (MAXISCQTDATA[207], MAXISCQTDATA_OUT[207]);
  buf B_MAXISCQTDATA208 (MAXISCQTDATA[208], MAXISCQTDATA_OUT[208]);
  buf B_MAXISCQTDATA209 (MAXISCQTDATA[209], MAXISCQTDATA_OUT[209]);
  buf B_MAXISCQTDATA21 (MAXISCQTDATA[21], MAXISCQTDATA_OUT[21]);
  buf B_MAXISCQTDATA210 (MAXISCQTDATA[210], MAXISCQTDATA_OUT[210]);
  buf B_MAXISCQTDATA211 (MAXISCQTDATA[211], MAXISCQTDATA_OUT[211]);
  buf B_MAXISCQTDATA212 (MAXISCQTDATA[212], MAXISCQTDATA_OUT[212]);
  buf B_MAXISCQTDATA213 (MAXISCQTDATA[213], MAXISCQTDATA_OUT[213]);
  buf B_MAXISCQTDATA214 (MAXISCQTDATA[214], MAXISCQTDATA_OUT[214]);
  buf B_MAXISCQTDATA215 (MAXISCQTDATA[215], MAXISCQTDATA_OUT[215]);
  buf B_MAXISCQTDATA216 (MAXISCQTDATA[216], MAXISCQTDATA_OUT[216]);
  buf B_MAXISCQTDATA217 (MAXISCQTDATA[217], MAXISCQTDATA_OUT[217]);
  buf B_MAXISCQTDATA218 (MAXISCQTDATA[218], MAXISCQTDATA_OUT[218]);
  buf B_MAXISCQTDATA219 (MAXISCQTDATA[219], MAXISCQTDATA_OUT[219]);
  buf B_MAXISCQTDATA22 (MAXISCQTDATA[22], MAXISCQTDATA_OUT[22]);
  buf B_MAXISCQTDATA220 (MAXISCQTDATA[220], MAXISCQTDATA_OUT[220]);
  buf B_MAXISCQTDATA221 (MAXISCQTDATA[221], MAXISCQTDATA_OUT[221]);
  buf B_MAXISCQTDATA222 (MAXISCQTDATA[222], MAXISCQTDATA_OUT[222]);
  buf B_MAXISCQTDATA223 (MAXISCQTDATA[223], MAXISCQTDATA_OUT[223]);
  buf B_MAXISCQTDATA224 (MAXISCQTDATA[224], MAXISCQTDATA_OUT[224]);
  buf B_MAXISCQTDATA225 (MAXISCQTDATA[225], MAXISCQTDATA_OUT[225]);
  buf B_MAXISCQTDATA226 (MAXISCQTDATA[226], MAXISCQTDATA_OUT[226]);
  buf B_MAXISCQTDATA227 (MAXISCQTDATA[227], MAXISCQTDATA_OUT[227]);
  buf B_MAXISCQTDATA228 (MAXISCQTDATA[228], MAXISCQTDATA_OUT[228]);
  buf B_MAXISCQTDATA229 (MAXISCQTDATA[229], MAXISCQTDATA_OUT[229]);
  buf B_MAXISCQTDATA23 (MAXISCQTDATA[23], MAXISCQTDATA_OUT[23]);
  buf B_MAXISCQTDATA230 (MAXISCQTDATA[230], MAXISCQTDATA_OUT[230]);
  buf B_MAXISCQTDATA231 (MAXISCQTDATA[231], MAXISCQTDATA_OUT[231]);
  buf B_MAXISCQTDATA232 (MAXISCQTDATA[232], MAXISCQTDATA_OUT[232]);
  buf B_MAXISCQTDATA233 (MAXISCQTDATA[233], MAXISCQTDATA_OUT[233]);
  buf B_MAXISCQTDATA234 (MAXISCQTDATA[234], MAXISCQTDATA_OUT[234]);
  buf B_MAXISCQTDATA235 (MAXISCQTDATA[235], MAXISCQTDATA_OUT[235]);
  buf B_MAXISCQTDATA236 (MAXISCQTDATA[236], MAXISCQTDATA_OUT[236]);
  buf B_MAXISCQTDATA237 (MAXISCQTDATA[237], MAXISCQTDATA_OUT[237]);
  buf B_MAXISCQTDATA238 (MAXISCQTDATA[238], MAXISCQTDATA_OUT[238]);
  buf B_MAXISCQTDATA239 (MAXISCQTDATA[239], MAXISCQTDATA_OUT[239]);
  buf B_MAXISCQTDATA24 (MAXISCQTDATA[24], MAXISCQTDATA_OUT[24]);
  buf B_MAXISCQTDATA240 (MAXISCQTDATA[240], MAXISCQTDATA_OUT[240]);
  buf B_MAXISCQTDATA241 (MAXISCQTDATA[241], MAXISCQTDATA_OUT[241]);
  buf B_MAXISCQTDATA242 (MAXISCQTDATA[242], MAXISCQTDATA_OUT[242]);
  buf B_MAXISCQTDATA243 (MAXISCQTDATA[243], MAXISCQTDATA_OUT[243]);
  buf B_MAXISCQTDATA244 (MAXISCQTDATA[244], MAXISCQTDATA_OUT[244]);
  buf B_MAXISCQTDATA245 (MAXISCQTDATA[245], MAXISCQTDATA_OUT[245]);
  buf B_MAXISCQTDATA246 (MAXISCQTDATA[246], MAXISCQTDATA_OUT[246]);
  buf B_MAXISCQTDATA247 (MAXISCQTDATA[247], MAXISCQTDATA_OUT[247]);
  buf B_MAXISCQTDATA248 (MAXISCQTDATA[248], MAXISCQTDATA_OUT[248]);
  buf B_MAXISCQTDATA249 (MAXISCQTDATA[249], MAXISCQTDATA_OUT[249]);
  buf B_MAXISCQTDATA25 (MAXISCQTDATA[25], MAXISCQTDATA_OUT[25]);
  buf B_MAXISCQTDATA250 (MAXISCQTDATA[250], MAXISCQTDATA_OUT[250]);
  buf B_MAXISCQTDATA251 (MAXISCQTDATA[251], MAXISCQTDATA_OUT[251]);
  buf B_MAXISCQTDATA252 (MAXISCQTDATA[252], MAXISCQTDATA_OUT[252]);
  buf B_MAXISCQTDATA253 (MAXISCQTDATA[253], MAXISCQTDATA_OUT[253]);
  buf B_MAXISCQTDATA254 (MAXISCQTDATA[254], MAXISCQTDATA_OUT[254]);
  buf B_MAXISCQTDATA255 (MAXISCQTDATA[255], MAXISCQTDATA_OUT[255]);
  buf B_MAXISCQTDATA26 (MAXISCQTDATA[26], MAXISCQTDATA_OUT[26]);
  buf B_MAXISCQTDATA27 (MAXISCQTDATA[27], MAXISCQTDATA_OUT[27]);
  buf B_MAXISCQTDATA28 (MAXISCQTDATA[28], MAXISCQTDATA_OUT[28]);
  buf B_MAXISCQTDATA29 (MAXISCQTDATA[29], MAXISCQTDATA_OUT[29]);
  buf B_MAXISCQTDATA3 (MAXISCQTDATA[3], MAXISCQTDATA_OUT[3]);
  buf B_MAXISCQTDATA30 (MAXISCQTDATA[30], MAXISCQTDATA_OUT[30]);
  buf B_MAXISCQTDATA31 (MAXISCQTDATA[31], MAXISCQTDATA_OUT[31]);
  buf B_MAXISCQTDATA32 (MAXISCQTDATA[32], MAXISCQTDATA_OUT[32]);
  buf B_MAXISCQTDATA33 (MAXISCQTDATA[33], MAXISCQTDATA_OUT[33]);
  buf B_MAXISCQTDATA34 (MAXISCQTDATA[34], MAXISCQTDATA_OUT[34]);
  buf B_MAXISCQTDATA35 (MAXISCQTDATA[35], MAXISCQTDATA_OUT[35]);
  buf B_MAXISCQTDATA36 (MAXISCQTDATA[36], MAXISCQTDATA_OUT[36]);
  buf B_MAXISCQTDATA37 (MAXISCQTDATA[37], MAXISCQTDATA_OUT[37]);
  buf B_MAXISCQTDATA38 (MAXISCQTDATA[38], MAXISCQTDATA_OUT[38]);
  buf B_MAXISCQTDATA39 (MAXISCQTDATA[39], MAXISCQTDATA_OUT[39]);
  buf B_MAXISCQTDATA4 (MAXISCQTDATA[4], MAXISCQTDATA_OUT[4]);
  buf B_MAXISCQTDATA40 (MAXISCQTDATA[40], MAXISCQTDATA_OUT[40]);
  buf B_MAXISCQTDATA41 (MAXISCQTDATA[41], MAXISCQTDATA_OUT[41]);
  buf B_MAXISCQTDATA42 (MAXISCQTDATA[42], MAXISCQTDATA_OUT[42]);
  buf B_MAXISCQTDATA43 (MAXISCQTDATA[43], MAXISCQTDATA_OUT[43]);
  buf B_MAXISCQTDATA44 (MAXISCQTDATA[44], MAXISCQTDATA_OUT[44]);
  buf B_MAXISCQTDATA45 (MAXISCQTDATA[45], MAXISCQTDATA_OUT[45]);
  buf B_MAXISCQTDATA46 (MAXISCQTDATA[46], MAXISCQTDATA_OUT[46]);
  buf B_MAXISCQTDATA47 (MAXISCQTDATA[47], MAXISCQTDATA_OUT[47]);
  buf B_MAXISCQTDATA48 (MAXISCQTDATA[48], MAXISCQTDATA_OUT[48]);
  buf B_MAXISCQTDATA49 (MAXISCQTDATA[49], MAXISCQTDATA_OUT[49]);
  buf B_MAXISCQTDATA5 (MAXISCQTDATA[5], MAXISCQTDATA_OUT[5]);
  buf B_MAXISCQTDATA50 (MAXISCQTDATA[50], MAXISCQTDATA_OUT[50]);
  buf B_MAXISCQTDATA51 (MAXISCQTDATA[51], MAXISCQTDATA_OUT[51]);
  buf B_MAXISCQTDATA52 (MAXISCQTDATA[52], MAXISCQTDATA_OUT[52]);
  buf B_MAXISCQTDATA53 (MAXISCQTDATA[53], MAXISCQTDATA_OUT[53]);
  buf B_MAXISCQTDATA54 (MAXISCQTDATA[54], MAXISCQTDATA_OUT[54]);
  buf B_MAXISCQTDATA55 (MAXISCQTDATA[55], MAXISCQTDATA_OUT[55]);
  buf B_MAXISCQTDATA56 (MAXISCQTDATA[56], MAXISCQTDATA_OUT[56]);
  buf B_MAXISCQTDATA57 (MAXISCQTDATA[57], MAXISCQTDATA_OUT[57]);
  buf B_MAXISCQTDATA58 (MAXISCQTDATA[58], MAXISCQTDATA_OUT[58]);
  buf B_MAXISCQTDATA59 (MAXISCQTDATA[59], MAXISCQTDATA_OUT[59]);
  buf B_MAXISCQTDATA6 (MAXISCQTDATA[6], MAXISCQTDATA_OUT[6]);
  buf B_MAXISCQTDATA60 (MAXISCQTDATA[60], MAXISCQTDATA_OUT[60]);
  buf B_MAXISCQTDATA61 (MAXISCQTDATA[61], MAXISCQTDATA_OUT[61]);
  buf B_MAXISCQTDATA62 (MAXISCQTDATA[62], MAXISCQTDATA_OUT[62]);
  buf B_MAXISCQTDATA63 (MAXISCQTDATA[63], MAXISCQTDATA_OUT[63]);
  buf B_MAXISCQTDATA64 (MAXISCQTDATA[64], MAXISCQTDATA_OUT[64]);
  buf B_MAXISCQTDATA65 (MAXISCQTDATA[65], MAXISCQTDATA_OUT[65]);
  buf B_MAXISCQTDATA66 (MAXISCQTDATA[66], MAXISCQTDATA_OUT[66]);
  buf B_MAXISCQTDATA67 (MAXISCQTDATA[67], MAXISCQTDATA_OUT[67]);
  buf B_MAXISCQTDATA68 (MAXISCQTDATA[68], MAXISCQTDATA_OUT[68]);
  buf B_MAXISCQTDATA69 (MAXISCQTDATA[69], MAXISCQTDATA_OUT[69]);
  buf B_MAXISCQTDATA7 (MAXISCQTDATA[7], MAXISCQTDATA_OUT[7]);
  buf B_MAXISCQTDATA70 (MAXISCQTDATA[70], MAXISCQTDATA_OUT[70]);
  buf B_MAXISCQTDATA71 (MAXISCQTDATA[71], MAXISCQTDATA_OUT[71]);
  buf B_MAXISCQTDATA72 (MAXISCQTDATA[72], MAXISCQTDATA_OUT[72]);
  buf B_MAXISCQTDATA73 (MAXISCQTDATA[73], MAXISCQTDATA_OUT[73]);
  buf B_MAXISCQTDATA74 (MAXISCQTDATA[74], MAXISCQTDATA_OUT[74]);
  buf B_MAXISCQTDATA75 (MAXISCQTDATA[75], MAXISCQTDATA_OUT[75]);
  buf B_MAXISCQTDATA76 (MAXISCQTDATA[76], MAXISCQTDATA_OUT[76]);
  buf B_MAXISCQTDATA77 (MAXISCQTDATA[77], MAXISCQTDATA_OUT[77]);
  buf B_MAXISCQTDATA78 (MAXISCQTDATA[78], MAXISCQTDATA_OUT[78]);
  buf B_MAXISCQTDATA79 (MAXISCQTDATA[79], MAXISCQTDATA_OUT[79]);
  buf B_MAXISCQTDATA8 (MAXISCQTDATA[8], MAXISCQTDATA_OUT[8]);
  buf B_MAXISCQTDATA80 (MAXISCQTDATA[80], MAXISCQTDATA_OUT[80]);
  buf B_MAXISCQTDATA81 (MAXISCQTDATA[81], MAXISCQTDATA_OUT[81]);
  buf B_MAXISCQTDATA82 (MAXISCQTDATA[82], MAXISCQTDATA_OUT[82]);
  buf B_MAXISCQTDATA83 (MAXISCQTDATA[83], MAXISCQTDATA_OUT[83]);
  buf B_MAXISCQTDATA84 (MAXISCQTDATA[84], MAXISCQTDATA_OUT[84]);
  buf B_MAXISCQTDATA85 (MAXISCQTDATA[85], MAXISCQTDATA_OUT[85]);
  buf B_MAXISCQTDATA86 (MAXISCQTDATA[86], MAXISCQTDATA_OUT[86]);
  buf B_MAXISCQTDATA87 (MAXISCQTDATA[87], MAXISCQTDATA_OUT[87]);
  buf B_MAXISCQTDATA88 (MAXISCQTDATA[88], MAXISCQTDATA_OUT[88]);
  buf B_MAXISCQTDATA89 (MAXISCQTDATA[89], MAXISCQTDATA_OUT[89]);
  buf B_MAXISCQTDATA9 (MAXISCQTDATA[9], MAXISCQTDATA_OUT[9]);
  buf B_MAXISCQTDATA90 (MAXISCQTDATA[90], MAXISCQTDATA_OUT[90]);
  buf B_MAXISCQTDATA91 (MAXISCQTDATA[91], MAXISCQTDATA_OUT[91]);
  buf B_MAXISCQTDATA92 (MAXISCQTDATA[92], MAXISCQTDATA_OUT[92]);
  buf B_MAXISCQTDATA93 (MAXISCQTDATA[93], MAXISCQTDATA_OUT[93]);
  buf B_MAXISCQTDATA94 (MAXISCQTDATA[94], MAXISCQTDATA_OUT[94]);
  buf B_MAXISCQTDATA95 (MAXISCQTDATA[95], MAXISCQTDATA_OUT[95]);
  buf B_MAXISCQTDATA96 (MAXISCQTDATA[96], MAXISCQTDATA_OUT[96]);
  buf B_MAXISCQTDATA97 (MAXISCQTDATA[97], MAXISCQTDATA_OUT[97]);
  buf B_MAXISCQTDATA98 (MAXISCQTDATA[98], MAXISCQTDATA_OUT[98]);
  buf B_MAXISCQTDATA99 (MAXISCQTDATA[99], MAXISCQTDATA_OUT[99]);
  buf B_MAXISCQTKEEP0 (MAXISCQTKEEP[0], MAXISCQTKEEP_OUT[0]);
  buf B_MAXISCQTKEEP1 (MAXISCQTKEEP[1], MAXISCQTKEEP_OUT[1]);
  buf B_MAXISCQTKEEP2 (MAXISCQTKEEP[2], MAXISCQTKEEP_OUT[2]);
  buf B_MAXISCQTKEEP3 (MAXISCQTKEEP[3], MAXISCQTKEEP_OUT[3]);
  buf B_MAXISCQTKEEP4 (MAXISCQTKEEP[4], MAXISCQTKEEP_OUT[4]);
  buf B_MAXISCQTKEEP5 (MAXISCQTKEEP[5], MAXISCQTKEEP_OUT[5]);
  buf B_MAXISCQTKEEP6 (MAXISCQTKEEP[6], MAXISCQTKEEP_OUT[6]);
  buf B_MAXISCQTKEEP7 (MAXISCQTKEEP[7], MAXISCQTKEEP_OUT[7]);
  buf B_MAXISCQTLAST (MAXISCQTLAST, MAXISCQTLAST_OUT);
  buf B_MAXISCQTUSER0 (MAXISCQTUSER[0], MAXISCQTUSER_OUT[0]);
  buf B_MAXISCQTUSER1 (MAXISCQTUSER[1], MAXISCQTUSER_OUT[1]);
  buf B_MAXISCQTUSER10 (MAXISCQTUSER[10], MAXISCQTUSER_OUT[10]);
  buf B_MAXISCQTUSER11 (MAXISCQTUSER[11], MAXISCQTUSER_OUT[11]);
  buf B_MAXISCQTUSER12 (MAXISCQTUSER[12], MAXISCQTUSER_OUT[12]);
  buf B_MAXISCQTUSER13 (MAXISCQTUSER[13], MAXISCQTUSER_OUT[13]);
  buf B_MAXISCQTUSER14 (MAXISCQTUSER[14], MAXISCQTUSER_OUT[14]);
  buf B_MAXISCQTUSER15 (MAXISCQTUSER[15], MAXISCQTUSER_OUT[15]);
  buf B_MAXISCQTUSER16 (MAXISCQTUSER[16], MAXISCQTUSER_OUT[16]);
  buf B_MAXISCQTUSER17 (MAXISCQTUSER[17], MAXISCQTUSER_OUT[17]);
  buf B_MAXISCQTUSER18 (MAXISCQTUSER[18], MAXISCQTUSER_OUT[18]);
  buf B_MAXISCQTUSER19 (MAXISCQTUSER[19], MAXISCQTUSER_OUT[19]);
  buf B_MAXISCQTUSER2 (MAXISCQTUSER[2], MAXISCQTUSER_OUT[2]);
  buf B_MAXISCQTUSER20 (MAXISCQTUSER[20], MAXISCQTUSER_OUT[20]);
  buf B_MAXISCQTUSER21 (MAXISCQTUSER[21], MAXISCQTUSER_OUT[21]);
  buf B_MAXISCQTUSER22 (MAXISCQTUSER[22], MAXISCQTUSER_OUT[22]);
  buf B_MAXISCQTUSER23 (MAXISCQTUSER[23], MAXISCQTUSER_OUT[23]);
  buf B_MAXISCQTUSER24 (MAXISCQTUSER[24], MAXISCQTUSER_OUT[24]);
  buf B_MAXISCQTUSER25 (MAXISCQTUSER[25], MAXISCQTUSER_OUT[25]);
  buf B_MAXISCQTUSER26 (MAXISCQTUSER[26], MAXISCQTUSER_OUT[26]);
  buf B_MAXISCQTUSER27 (MAXISCQTUSER[27], MAXISCQTUSER_OUT[27]);
  buf B_MAXISCQTUSER28 (MAXISCQTUSER[28], MAXISCQTUSER_OUT[28]);
  buf B_MAXISCQTUSER29 (MAXISCQTUSER[29], MAXISCQTUSER_OUT[29]);
  buf B_MAXISCQTUSER3 (MAXISCQTUSER[3], MAXISCQTUSER_OUT[3]);
  buf B_MAXISCQTUSER30 (MAXISCQTUSER[30], MAXISCQTUSER_OUT[30]);
  buf B_MAXISCQTUSER31 (MAXISCQTUSER[31], MAXISCQTUSER_OUT[31]);
  buf B_MAXISCQTUSER32 (MAXISCQTUSER[32], MAXISCQTUSER_OUT[32]);
  buf B_MAXISCQTUSER33 (MAXISCQTUSER[33], MAXISCQTUSER_OUT[33]);
  buf B_MAXISCQTUSER34 (MAXISCQTUSER[34], MAXISCQTUSER_OUT[34]);
  buf B_MAXISCQTUSER35 (MAXISCQTUSER[35], MAXISCQTUSER_OUT[35]);
  buf B_MAXISCQTUSER36 (MAXISCQTUSER[36], MAXISCQTUSER_OUT[36]);
  buf B_MAXISCQTUSER37 (MAXISCQTUSER[37], MAXISCQTUSER_OUT[37]);
  buf B_MAXISCQTUSER38 (MAXISCQTUSER[38], MAXISCQTUSER_OUT[38]);
  buf B_MAXISCQTUSER39 (MAXISCQTUSER[39], MAXISCQTUSER_OUT[39]);
  buf B_MAXISCQTUSER4 (MAXISCQTUSER[4], MAXISCQTUSER_OUT[4]);
  buf B_MAXISCQTUSER40 (MAXISCQTUSER[40], MAXISCQTUSER_OUT[40]);
  buf B_MAXISCQTUSER41 (MAXISCQTUSER[41], MAXISCQTUSER_OUT[41]);
  buf B_MAXISCQTUSER42 (MAXISCQTUSER[42], MAXISCQTUSER_OUT[42]);
  buf B_MAXISCQTUSER43 (MAXISCQTUSER[43], MAXISCQTUSER_OUT[43]);
  buf B_MAXISCQTUSER44 (MAXISCQTUSER[44], MAXISCQTUSER_OUT[44]);
  buf B_MAXISCQTUSER45 (MAXISCQTUSER[45], MAXISCQTUSER_OUT[45]);
  buf B_MAXISCQTUSER46 (MAXISCQTUSER[46], MAXISCQTUSER_OUT[46]);
  buf B_MAXISCQTUSER47 (MAXISCQTUSER[47], MAXISCQTUSER_OUT[47]);
  buf B_MAXISCQTUSER48 (MAXISCQTUSER[48], MAXISCQTUSER_OUT[48]);
  buf B_MAXISCQTUSER49 (MAXISCQTUSER[49], MAXISCQTUSER_OUT[49]);
  buf B_MAXISCQTUSER5 (MAXISCQTUSER[5], MAXISCQTUSER_OUT[5]);
  buf B_MAXISCQTUSER50 (MAXISCQTUSER[50], MAXISCQTUSER_OUT[50]);
  buf B_MAXISCQTUSER51 (MAXISCQTUSER[51], MAXISCQTUSER_OUT[51]);
  buf B_MAXISCQTUSER52 (MAXISCQTUSER[52], MAXISCQTUSER_OUT[52]);
  buf B_MAXISCQTUSER53 (MAXISCQTUSER[53], MAXISCQTUSER_OUT[53]);
  buf B_MAXISCQTUSER54 (MAXISCQTUSER[54], MAXISCQTUSER_OUT[54]);
  buf B_MAXISCQTUSER55 (MAXISCQTUSER[55], MAXISCQTUSER_OUT[55]);
  buf B_MAXISCQTUSER56 (MAXISCQTUSER[56], MAXISCQTUSER_OUT[56]);
  buf B_MAXISCQTUSER57 (MAXISCQTUSER[57], MAXISCQTUSER_OUT[57]);
  buf B_MAXISCQTUSER58 (MAXISCQTUSER[58], MAXISCQTUSER_OUT[58]);
  buf B_MAXISCQTUSER59 (MAXISCQTUSER[59], MAXISCQTUSER_OUT[59]);
  buf B_MAXISCQTUSER6 (MAXISCQTUSER[6], MAXISCQTUSER_OUT[6]);
  buf B_MAXISCQTUSER60 (MAXISCQTUSER[60], MAXISCQTUSER_OUT[60]);
  buf B_MAXISCQTUSER61 (MAXISCQTUSER[61], MAXISCQTUSER_OUT[61]);
  buf B_MAXISCQTUSER62 (MAXISCQTUSER[62], MAXISCQTUSER_OUT[62]);
  buf B_MAXISCQTUSER63 (MAXISCQTUSER[63], MAXISCQTUSER_OUT[63]);
  buf B_MAXISCQTUSER64 (MAXISCQTUSER[64], MAXISCQTUSER_OUT[64]);
  buf B_MAXISCQTUSER65 (MAXISCQTUSER[65], MAXISCQTUSER_OUT[65]);
  buf B_MAXISCQTUSER66 (MAXISCQTUSER[66], MAXISCQTUSER_OUT[66]);
  buf B_MAXISCQTUSER67 (MAXISCQTUSER[67], MAXISCQTUSER_OUT[67]);
  buf B_MAXISCQTUSER68 (MAXISCQTUSER[68], MAXISCQTUSER_OUT[68]);
  buf B_MAXISCQTUSER69 (MAXISCQTUSER[69], MAXISCQTUSER_OUT[69]);
  buf B_MAXISCQTUSER7 (MAXISCQTUSER[7], MAXISCQTUSER_OUT[7]);
  buf B_MAXISCQTUSER70 (MAXISCQTUSER[70], MAXISCQTUSER_OUT[70]);
  buf B_MAXISCQTUSER71 (MAXISCQTUSER[71], MAXISCQTUSER_OUT[71]);
  buf B_MAXISCQTUSER72 (MAXISCQTUSER[72], MAXISCQTUSER_OUT[72]);
  buf B_MAXISCQTUSER73 (MAXISCQTUSER[73], MAXISCQTUSER_OUT[73]);
  buf B_MAXISCQTUSER74 (MAXISCQTUSER[74], MAXISCQTUSER_OUT[74]);
  buf B_MAXISCQTUSER75 (MAXISCQTUSER[75], MAXISCQTUSER_OUT[75]);
  buf B_MAXISCQTUSER76 (MAXISCQTUSER[76], MAXISCQTUSER_OUT[76]);
  buf B_MAXISCQTUSER77 (MAXISCQTUSER[77], MAXISCQTUSER_OUT[77]);
  buf B_MAXISCQTUSER78 (MAXISCQTUSER[78], MAXISCQTUSER_OUT[78]);
  buf B_MAXISCQTUSER79 (MAXISCQTUSER[79], MAXISCQTUSER_OUT[79]);
  buf B_MAXISCQTUSER8 (MAXISCQTUSER[8], MAXISCQTUSER_OUT[8]);
  buf B_MAXISCQTUSER80 (MAXISCQTUSER[80], MAXISCQTUSER_OUT[80]);
  buf B_MAXISCQTUSER81 (MAXISCQTUSER[81], MAXISCQTUSER_OUT[81]);
  buf B_MAXISCQTUSER82 (MAXISCQTUSER[82], MAXISCQTUSER_OUT[82]);
  buf B_MAXISCQTUSER83 (MAXISCQTUSER[83], MAXISCQTUSER_OUT[83]);
  buf B_MAXISCQTUSER84 (MAXISCQTUSER[84], MAXISCQTUSER_OUT[84]);
  buf B_MAXISCQTUSER9 (MAXISCQTUSER[9], MAXISCQTUSER_OUT[9]);
  buf B_MAXISCQTVALID (MAXISCQTVALID, MAXISCQTVALID_OUT);
  buf B_MAXISRCTDATA0 (MAXISRCTDATA[0], MAXISRCTDATA_OUT[0]);
  buf B_MAXISRCTDATA1 (MAXISRCTDATA[1], MAXISRCTDATA_OUT[1]);
  buf B_MAXISRCTDATA10 (MAXISRCTDATA[10], MAXISRCTDATA_OUT[10]);
  buf B_MAXISRCTDATA100 (MAXISRCTDATA[100], MAXISRCTDATA_OUT[100]);
  buf B_MAXISRCTDATA101 (MAXISRCTDATA[101], MAXISRCTDATA_OUT[101]);
  buf B_MAXISRCTDATA102 (MAXISRCTDATA[102], MAXISRCTDATA_OUT[102]);
  buf B_MAXISRCTDATA103 (MAXISRCTDATA[103], MAXISRCTDATA_OUT[103]);
  buf B_MAXISRCTDATA104 (MAXISRCTDATA[104], MAXISRCTDATA_OUT[104]);
  buf B_MAXISRCTDATA105 (MAXISRCTDATA[105], MAXISRCTDATA_OUT[105]);
  buf B_MAXISRCTDATA106 (MAXISRCTDATA[106], MAXISRCTDATA_OUT[106]);
  buf B_MAXISRCTDATA107 (MAXISRCTDATA[107], MAXISRCTDATA_OUT[107]);
  buf B_MAXISRCTDATA108 (MAXISRCTDATA[108], MAXISRCTDATA_OUT[108]);
  buf B_MAXISRCTDATA109 (MAXISRCTDATA[109], MAXISRCTDATA_OUT[109]);
  buf B_MAXISRCTDATA11 (MAXISRCTDATA[11], MAXISRCTDATA_OUT[11]);
  buf B_MAXISRCTDATA110 (MAXISRCTDATA[110], MAXISRCTDATA_OUT[110]);
  buf B_MAXISRCTDATA111 (MAXISRCTDATA[111], MAXISRCTDATA_OUT[111]);
  buf B_MAXISRCTDATA112 (MAXISRCTDATA[112], MAXISRCTDATA_OUT[112]);
  buf B_MAXISRCTDATA113 (MAXISRCTDATA[113], MAXISRCTDATA_OUT[113]);
  buf B_MAXISRCTDATA114 (MAXISRCTDATA[114], MAXISRCTDATA_OUT[114]);
  buf B_MAXISRCTDATA115 (MAXISRCTDATA[115], MAXISRCTDATA_OUT[115]);
  buf B_MAXISRCTDATA116 (MAXISRCTDATA[116], MAXISRCTDATA_OUT[116]);
  buf B_MAXISRCTDATA117 (MAXISRCTDATA[117], MAXISRCTDATA_OUT[117]);
  buf B_MAXISRCTDATA118 (MAXISRCTDATA[118], MAXISRCTDATA_OUT[118]);
  buf B_MAXISRCTDATA119 (MAXISRCTDATA[119], MAXISRCTDATA_OUT[119]);
  buf B_MAXISRCTDATA12 (MAXISRCTDATA[12], MAXISRCTDATA_OUT[12]);
  buf B_MAXISRCTDATA120 (MAXISRCTDATA[120], MAXISRCTDATA_OUT[120]);
  buf B_MAXISRCTDATA121 (MAXISRCTDATA[121], MAXISRCTDATA_OUT[121]);
  buf B_MAXISRCTDATA122 (MAXISRCTDATA[122], MAXISRCTDATA_OUT[122]);
  buf B_MAXISRCTDATA123 (MAXISRCTDATA[123], MAXISRCTDATA_OUT[123]);
  buf B_MAXISRCTDATA124 (MAXISRCTDATA[124], MAXISRCTDATA_OUT[124]);
  buf B_MAXISRCTDATA125 (MAXISRCTDATA[125], MAXISRCTDATA_OUT[125]);
  buf B_MAXISRCTDATA126 (MAXISRCTDATA[126], MAXISRCTDATA_OUT[126]);
  buf B_MAXISRCTDATA127 (MAXISRCTDATA[127], MAXISRCTDATA_OUT[127]);
  buf B_MAXISRCTDATA128 (MAXISRCTDATA[128], MAXISRCTDATA_OUT[128]);
  buf B_MAXISRCTDATA129 (MAXISRCTDATA[129], MAXISRCTDATA_OUT[129]);
  buf B_MAXISRCTDATA13 (MAXISRCTDATA[13], MAXISRCTDATA_OUT[13]);
  buf B_MAXISRCTDATA130 (MAXISRCTDATA[130], MAXISRCTDATA_OUT[130]);
  buf B_MAXISRCTDATA131 (MAXISRCTDATA[131], MAXISRCTDATA_OUT[131]);
  buf B_MAXISRCTDATA132 (MAXISRCTDATA[132], MAXISRCTDATA_OUT[132]);
  buf B_MAXISRCTDATA133 (MAXISRCTDATA[133], MAXISRCTDATA_OUT[133]);
  buf B_MAXISRCTDATA134 (MAXISRCTDATA[134], MAXISRCTDATA_OUT[134]);
  buf B_MAXISRCTDATA135 (MAXISRCTDATA[135], MAXISRCTDATA_OUT[135]);
  buf B_MAXISRCTDATA136 (MAXISRCTDATA[136], MAXISRCTDATA_OUT[136]);
  buf B_MAXISRCTDATA137 (MAXISRCTDATA[137], MAXISRCTDATA_OUT[137]);
  buf B_MAXISRCTDATA138 (MAXISRCTDATA[138], MAXISRCTDATA_OUT[138]);
  buf B_MAXISRCTDATA139 (MAXISRCTDATA[139], MAXISRCTDATA_OUT[139]);
  buf B_MAXISRCTDATA14 (MAXISRCTDATA[14], MAXISRCTDATA_OUT[14]);
  buf B_MAXISRCTDATA140 (MAXISRCTDATA[140], MAXISRCTDATA_OUT[140]);
  buf B_MAXISRCTDATA141 (MAXISRCTDATA[141], MAXISRCTDATA_OUT[141]);
  buf B_MAXISRCTDATA142 (MAXISRCTDATA[142], MAXISRCTDATA_OUT[142]);
  buf B_MAXISRCTDATA143 (MAXISRCTDATA[143], MAXISRCTDATA_OUT[143]);
  buf B_MAXISRCTDATA144 (MAXISRCTDATA[144], MAXISRCTDATA_OUT[144]);
  buf B_MAXISRCTDATA145 (MAXISRCTDATA[145], MAXISRCTDATA_OUT[145]);
  buf B_MAXISRCTDATA146 (MAXISRCTDATA[146], MAXISRCTDATA_OUT[146]);
  buf B_MAXISRCTDATA147 (MAXISRCTDATA[147], MAXISRCTDATA_OUT[147]);
  buf B_MAXISRCTDATA148 (MAXISRCTDATA[148], MAXISRCTDATA_OUT[148]);
  buf B_MAXISRCTDATA149 (MAXISRCTDATA[149], MAXISRCTDATA_OUT[149]);
  buf B_MAXISRCTDATA15 (MAXISRCTDATA[15], MAXISRCTDATA_OUT[15]);
  buf B_MAXISRCTDATA150 (MAXISRCTDATA[150], MAXISRCTDATA_OUT[150]);
  buf B_MAXISRCTDATA151 (MAXISRCTDATA[151], MAXISRCTDATA_OUT[151]);
  buf B_MAXISRCTDATA152 (MAXISRCTDATA[152], MAXISRCTDATA_OUT[152]);
  buf B_MAXISRCTDATA153 (MAXISRCTDATA[153], MAXISRCTDATA_OUT[153]);
  buf B_MAXISRCTDATA154 (MAXISRCTDATA[154], MAXISRCTDATA_OUT[154]);
  buf B_MAXISRCTDATA155 (MAXISRCTDATA[155], MAXISRCTDATA_OUT[155]);
  buf B_MAXISRCTDATA156 (MAXISRCTDATA[156], MAXISRCTDATA_OUT[156]);
  buf B_MAXISRCTDATA157 (MAXISRCTDATA[157], MAXISRCTDATA_OUT[157]);
  buf B_MAXISRCTDATA158 (MAXISRCTDATA[158], MAXISRCTDATA_OUT[158]);
  buf B_MAXISRCTDATA159 (MAXISRCTDATA[159], MAXISRCTDATA_OUT[159]);
  buf B_MAXISRCTDATA16 (MAXISRCTDATA[16], MAXISRCTDATA_OUT[16]);
  buf B_MAXISRCTDATA160 (MAXISRCTDATA[160], MAXISRCTDATA_OUT[160]);
  buf B_MAXISRCTDATA161 (MAXISRCTDATA[161], MAXISRCTDATA_OUT[161]);
  buf B_MAXISRCTDATA162 (MAXISRCTDATA[162], MAXISRCTDATA_OUT[162]);
  buf B_MAXISRCTDATA163 (MAXISRCTDATA[163], MAXISRCTDATA_OUT[163]);
  buf B_MAXISRCTDATA164 (MAXISRCTDATA[164], MAXISRCTDATA_OUT[164]);
  buf B_MAXISRCTDATA165 (MAXISRCTDATA[165], MAXISRCTDATA_OUT[165]);
  buf B_MAXISRCTDATA166 (MAXISRCTDATA[166], MAXISRCTDATA_OUT[166]);
  buf B_MAXISRCTDATA167 (MAXISRCTDATA[167], MAXISRCTDATA_OUT[167]);
  buf B_MAXISRCTDATA168 (MAXISRCTDATA[168], MAXISRCTDATA_OUT[168]);
  buf B_MAXISRCTDATA169 (MAXISRCTDATA[169], MAXISRCTDATA_OUT[169]);
  buf B_MAXISRCTDATA17 (MAXISRCTDATA[17], MAXISRCTDATA_OUT[17]);
  buf B_MAXISRCTDATA170 (MAXISRCTDATA[170], MAXISRCTDATA_OUT[170]);
  buf B_MAXISRCTDATA171 (MAXISRCTDATA[171], MAXISRCTDATA_OUT[171]);
  buf B_MAXISRCTDATA172 (MAXISRCTDATA[172], MAXISRCTDATA_OUT[172]);
  buf B_MAXISRCTDATA173 (MAXISRCTDATA[173], MAXISRCTDATA_OUT[173]);
  buf B_MAXISRCTDATA174 (MAXISRCTDATA[174], MAXISRCTDATA_OUT[174]);
  buf B_MAXISRCTDATA175 (MAXISRCTDATA[175], MAXISRCTDATA_OUT[175]);
  buf B_MAXISRCTDATA176 (MAXISRCTDATA[176], MAXISRCTDATA_OUT[176]);
  buf B_MAXISRCTDATA177 (MAXISRCTDATA[177], MAXISRCTDATA_OUT[177]);
  buf B_MAXISRCTDATA178 (MAXISRCTDATA[178], MAXISRCTDATA_OUT[178]);
  buf B_MAXISRCTDATA179 (MAXISRCTDATA[179], MAXISRCTDATA_OUT[179]);
  buf B_MAXISRCTDATA18 (MAXISRCTDATA[18], MAXISRCTDATA_OUT[18]);
  buf B_MAXISRCTDATA180 (MAXISRCTDATA[180], MAXISRCTDATA_OUT[180]);
  buf B_MAXISRCTDATA181 (MAXISRCTDATA[181], MAXISRCTDATA_OUT[181]);
  buf B_MAXISRCTDATA182 (MAXISRCTDATA[182], MAXISRCTDATA_OUT[182]);
  buf B_MAXISRCTDATA183 (MAXISRCTDATA[183], MAXISRCTDATA_OUT[183]);
  buf B_MAXISRCTDATA184 (MAXISRCTDATA[184], MAXISRCTDATA_OUT[184]);
  buf B_MAXISRCTDATA185 (MAXISRCTDATA[185], MAXISRCTDATA_OUT[185]);
  buf B_MAXISRCTDATA186 (MAXISRCTDATA[186], MAXISRCTDATA_OUT[186]);
  buf B_MAXISRCTDATA187 (MAXISRCTDATA[187], MAXISRCTDATA_OUT[187]);
  buf B_MAXISRCTDATA188 (MAXISRCTDATA[188], MAXISRCTDATA_OUT[188]);
  buf B_MAXISRCTDATA189 (MAXISRCTDATA[189], MAXISRCTDATA_OUT[189]);
  buf B_MAXISRCTDATA19 (MAXISRCTDATA[19], MAXISRCTDATA_OUT[19]);
  buf B_MAXISRCTDATA190 (MAXISRCTDATA[190], MAXISRCTDATA_OUT[190]);
  buf B_MAXISRCTDATA191 (MAXISRCTDATA[191], MAXISRCTDATA_OUT[191]);
  buf B_MAXISRCTDATA192 (MAXISRCTDATA[192], MAXISRCTDATA_OUT[192]);
  buf B_MAXISRCTDATA193 (MAXISRCTDATA[193], MAXISRCTDATA_OUT[193]);
  buf B_MAXISRCTDATA194 (MAXISRCTDATA[194], MAXISRCTDATA_OUT[194]);
  buf B_MAXISRCTDATA195 (MAXISRCTDATA[195], MAXISRCTDATA_OUT[195]);
  buf B_MAXISRCTDATA196 (MAXISRCTDATA[196], MAXISRCTDATA_OUT[196]);
  buf B_MAXISRCTDATA197 (MAXISRCTDATA[197], MAXISRCTDATA_OUT[197]);
  buf B_MAXISRCTDATA198 (MAXISRCTDATA[198], MAXISRCTDATA_OUT[198]);
  buf B_MAXISRCTDATA199 (MAXISRCTDATA[199], MAXISRCTDATA_OUT[199]);
  buf B_MAXISRCTDATA2 (MAXISRCTDATA[2], MAXISRCTDATA_OUT[2]);
  buf B_MAXISRCTDATA20 (MAXISRCTDATA[20], MAXISRCTDATA_OUT[20]);
  buf B_MAXISRCTDATA200 (MAXISRCTDATA[200], MAXISRCTDATA_OUT[200]);
  buf B_MAXISRCTDATA201 (MAXISRCTDATA[201], MAXISRCTDATA_OUT[201]);
  buf B_MAXISRCTDATA202 (MAXISRCTDATA[202], MAXISRCTDATA_OUT[202]);
  buf B_MAXISRCTDATA203 (MAXISRCTDATA[203], MAXISRCTDATA_OUT[203]);
  buf B_MAXISRCTDATA204 (MAXISRCTDATA[204], MAXISRCTDATA_OUT[204]);
  buf B_MAXISRCTDATA205 (MAXISRCTDATA[205], MAXISRCTDATA_OUT[205]);
  buf B_MAXISRCTDATA206 (MAXISRCTDATA[206], MAXISRCTDATA_OUT[206]);
  buf B_MAXISRCTDATA207 (MAXISRCTDATA[207], MAXISRCTDATA_OUT[207]);
  buf B_MAXISRCTDATA208 (MAXISRCTDATA[208], MAXISRCTDATA_OUT[208]);
  buf B_MAXISRCTDATA209 (MAXISRCTDATA[209], MAXISRCTDATA_OUT[209]);
  buf B_MAXISRCTDATA21 (MAXISRCTDATA[21], MAXISRCTDATA_OUT[21]);
  buf B_MAXISRCTDATA210 (MAXISRCTDATA[210], MAXISRCTDATA_OUT[210]);
  buf B_MAXISRCTDATA211 (MAXISRCTDATA[211], MAXISRCTDATA_OUT[211]);
  buf B_MAXISRCTDATA212 (MAXISRCTDATA[212], MAXISRCTDATA_OUT[212]);
  buf B_MAXISRCTDATA213 (MAXISRCTDATA[213], MAXISRCTDATA_OUT[213]);
  buf B_MAXISRCTDATA214 (MAXISRCTDATA[214], MAXISRCTDATA_OUT[214]);
  buf B_MAXISRCTDATA215 (MAXISRCTDATA[215], MAXISRCTDATA_OUT[215]);
  buf B_MAXISRCTDATA216 (MAXISRCTDATA[216], MAXISRCTDATA_OUT[216]);
  buf B_MAXISRCTDATA217 (MAXISRCTDATA[217], MAXISRCTDATA_OUT[217]);
  buf B_MAXISRCTDATA218 (MAXISRCTDATA[218], MAXISRCTDATA_OUT[218]);
  buf B_MAXISRCTDATA219 (MAXISRCTDATA[219], MAXISRCTDATA_OUT[219]);
  buf B_MAXISRCTDATA22 (MAXISRCTDATA[22], MAXISRCTDATA_OUT[22]);
  buf B_MAXISRCTDATA220 (MAXISRCTDATA[220], MAXISRCTDATA_OUT[220]);
  buf B_MAXISRCTDATA221 (MAXISRCTDATA[221], MAXISRCTDATA_OUT[221]);
  buf B_MAXISRCTDATA222 (MAXISRCTDATA[222], MAXISRCTDATA_OUT[222]);
  buf B_MAXISRCTDATA223 (MAXISRCTDATA[223], MAXISRCTDATA_OUT[223]);
  buf B_MAXISRCTDATA224 (MAXISRCTDATA[224], MAXISRCTDATA_OUT[224]);
  buf B_MAXISRCTDATA225 (MAXISRCTDATA[225], MAXISRCTDATA_OUT[225]);
  buf B_MAXISRCTDATA226 (MAXISRCTDATA[226], MAXISRCTDATA_OUT[226]);
  buf B_MAXISRCTDATA227 (MAXISRCTDATA[227], MAXISRCTDATA_OUT[227]);
  buf B_MAXISRCTDATA228 (MAXISRCTDATA[228], MAXISRCTDATA_OUT[228]);
  buf B_MAXISRCTDATA229 (MAXISRCTDATA[229], MAXISRCTDATA_OUT[229]);
  buf B_MAXISRCTDATA23 (MAXISRCTDATA[23], MAXISRCTDATA_OUT[23]);
  buf B_MAXISRCTDATA230 (MAXISRCTDATA[230], MAXISRCTDATA_OUT[230]);
  buf B_MAXISRCTDATA231 (MAXISRCTDATA[231], MAXISRCTDATA_OUT[231]);
  buf B_MAXISRCTDATA232 (MAXISRCTDATA[232], MAXISRCTDATA_OUT[232]);
  buf B_MAXISRCTDATA233 (MAXISRCTDATA[233], MAXISRCTDATA_OUT[233]);
  buf B_MAXISRCTDATA234 (MAXISRCTDATA[234], MAXISRCTDATA_OUT[234]);
  buf B_MAXISRCTDATA235 (MAXISRCTDATA[235], MAXISRCTDATA_OUT[235]);
  buf B_MAXISRCTDATA236 (MAXISRCTDATA[236], MAXISRCTDATA_OUT[236]);
  buf B_MAXISRCTDATA237 (MAXISRCTDATA[237], MAXISRCTDATA_OUT[237]);
  buf B_MAXISRCTDATA238 (MAXISRCTDATA[238], MAXISRCTDATA_OUT[238]);
  buf B_MAXISRCTDATA239 (MAXISRCTDATA[239], MAXISRCTDATA_OUT[239]);
  buf B_MAXISRCTDATA24 (MAXISRCTDATA[24], MAXISRCTDATA_OUT[24]);
  buf B_MAXISRCTDATA240 (MAXISRCTDATA[240], MAXISRCTDATA_OUT[240]);
  buf B_MAXISRCTDATA241 (MAXISRCTDATA[241], MAXISRCTDATA_OUT[241]);
  buf B_MAXISRCTDATA242 (MAXISRCTDATA[242], MAXISRCTDATA_OUT[242]);
  buf B_MAXISRCTDATA243 (MAXISRCTDATA[243], MAXISRCTDATA_OUT[243]);
  buf B_MAXISRCTDATA244 (MAXISRCTDATA[244], MAXISRCTDATA_OUT[244]);
  buf B_MAXISRCTDATA245 (MAXISRCTDATA[245], MAXISRCTDATA_OUT[245]);
  buf B_MAXISRCTDATA246 (MAXISRCTDATA[246], MAXISRCTDATA_OUT[246]);
  buf B_MAXISRCTDATA247 (MAXISRCTDATA[247], MAXISRCTDATA_OUT[247]);
  buf B_MAXISRCTDATA248 (MAXISRCTDATA[248], MAXISRCTDATA_OUT[248]);
  buf B_MAXISRCTDATA249 (MAXISRCTDATA[249], MAXISRCTDATA_OUT[249]);
  buf B_MAXISRCTDATA25 (MAXISRCTDATA[25], MAXISRCTDATA_OUT[25]);
  buf B_MAXISRCTDATA250 (MAXISRCTDATA[250], MAXISRCTDATA_OUT[250]);
  buf B_MAXISRCTDATA251 (MAXISRCTDATA[251], MAXISRCTDATA_OUT[251]);
  buf B_MAXISRCTDATA252 (MAXISRCTDATA[252], MAXISRCTDATA_OUT[252]);
  buf B_MAXISRCTDATA253 (MAXISRCTDATA[253], MAXISRCTDATA_OUT[253]);
  buf B_MAXISRCTDATA254 (MAXISRCTDATA[254], MAXISRCTDATA_OUT[254]);
  buf B_MAXISRCTDATA255 (MAXISRCTDATA[255], MAXISRCTDATA_OUT[255]);
  buf B_MAXISRCTDATA26 (MAXISRCTDATA[26], MAXISRCTDATA_OUT[26]);
  buf B_MAXISRCTDATA27 (MAXISRCTDATA[27], MAXISRCTDATA_OUT[27]);
  buf B_MAXISRCTDATA28 (MAXISRCTDATA[28], MAXISRCTDATA_OUT[28]);
  buf B_MAXISRCTDATA29 (MAXISRCTDATA[29], MAXISRCTDATA_OUT[29]);
  buf B_MAXISRCTDATA3 (MAXISRCTDATA[3], MAXISRCTDATA_OUT[3]);
  buf B_MAXISRCTDATA30 (MAXISRCTDATA[30], MAXISRCTDATA_OUT[30]);
  buf B_MAXISRCTDATA31 (MAXISRCTDATA[31], MAXISRCTDATA_OUT[31]);
  buf B_MAXISRCTDATA32 (MAXISRCTDATA[32], MAXISRCTDATA_OUT[32]);
  buf B_MAXISRCTDATA33 (MAXISRCTDATA[33], MAXISRCTDATA_OUT[33]);
  buf B_MAXISRCTDATA34 (MAXISRCTDATA[34], MAXISRCTDATA_OUT[34]);
  buf B_MAXISRCTDATA35 (MAXISRCTDATA[35], MAXISRCTDATA_OUT[35]);
  buf B_MAXISRCTDATA36 (MAXISRCTDATA[36], MAXISRCTDATA_OUT[36]);
  buf B_MAXISRCTDATA37 (MAXISRCTDATA[37], MAXISRCTDATA_OUT[37]);
  buf B_MAXISRCTDATA38 (MAXISRCTDATA[38], MAXISRCTDATA_OUT[38]);
  buf B_MAXISRCTDATA39 (MAXISRCTDATA[39], MAXISRCTDATA_OUT[39]);
  buf B_MAXISRCTDATA4 (MAXISRCTDATA[4], MAXISRCTDATA_OUT[4]);
  buf B_MAXISRCTDATA40 (MAXISRCTDATA[40], MAXISRCTDATA_OUT[40]);
  buf B_MAXISRCTDATA41 (MAXISRCTDATA[41], MAXISRCTDATA_OUT[41]);
  buf B_MAXISRCTDATA42 (MAXISRCTDATA[42], MAXISRCTDATA_OUT[42]);
  buf B_MAXISRCTDATA43 (MAXISRCTDATA[43], MAXISRCTDATA_OUT[43]);
  buf B_MAXISRCTDATA44 (MAXISRCTDATA[44], MAXISRCTDATA_OUT[44]);
  buf B_MAXISRCTDATA45 (MAXISRCTDATA[45], MAXISRCTDATA_OUT[45]);
  buf B_MAXISRCTDATA46 (MAXISRCTDATA[46], MAXISRCTDATA_OUT[46]);
  buf B_MAXISRCTDATA47 (MAXISRCTDATA[47], MAXISRCTDATA_OUT[47]);
  buf B_MAXISRCTDATA48 (MAXISRCTDATA[48], MAXISRCTDATA_OUT[48]);
  buf B_MAXISRCTDATA49 (MAXISRCTDATA[49], MAXISRCTDATA_OUT[49]);
  buf B_MAXISRCTDATA5 (MAXISRCTDATA[5], MAXISRCTDATA_OUT[5]);
  buf B_MAXISRCTDATA50 (MAXISRCTDATA[50], MAXISRCTDATA_OUT[50]);
  buf B_MAXISRCTDATA51 (MAXISRCTDATA[51], MAXISRCTDATA_OUT[51]);
  buf B_MAXISRCTDATA52 (MAXISRCTDATA[52], MAXISRCTDATA_OUT[52]);
  buf B_MAXISRCTDATA53 (MAXISRCTDATA[53], MAXISRCTDATA_OUT[53]);
  buf B_MAXISRCTDATA54 (MAXISRCTDATA[54], MAXISRCTDATA_OUT[54]);
  buf B_MAXISRCTDATA55 (MAXISRCTDATA[55], MAXISRCTDATA_OUT[55]);
  buf B_MAXISRCTDATA56 (MAXISRCTDATA[56], MAXISRCTDATA_OUT[56]);
  buf B_MAXISRCTDATA57 (MAXISRCTDATA[57], MAXISRCTDATA_OUT[57]);
  buf B_MAXISRCTDATA58 (MAXISRCTDATA[58], MAXISRCTDATA_OUT[58]);
  buf B_MAXISRCTDATA59 (MAXISRCTDATA[59], MAXISRCTDATA_OUT[59]);
  buf B_MAXISRCTDATA6 (MAXISRCTDATA[6], MAXISRCTDATA_OUT[6]);
  buf B_MAXISRCTDATA60 (MAXISRCTDATA[60], MAXISRCTDATA_OUT[60]);
  buf B_MAXISRCTDATA61 (MAXISRCTDATA[61], MAXISRCTDATA_OUT[61]);
  buf B_MAXISRCTDATA62 (MAXISRCTDATA[62], MAXISRCTDATA_OUT[62]);
  buf B_MAXISRCTDATA63 (MAXISRCTDATA[63], MAXISRCTDATA_OUT[63]);
  buf B_MAXISRCTDATA64 (MAXISRCTDATA[64], MAXISRCTDATA_OUT[64]);
  buf B_MAXISRCTDATA65 (MAXISRCTDATA[65], MAXISRCTDATA_OUT[65]);
  buf B_MAXISRCTDATA66 (MAXISRCTDATA[66], MAXISRCTDATA_OUT[66]);
  buf B_MAXISRCTDATA67 (MAXISRCTDATA[67], MAXISRCTDATA_OUT[67]);
  buf B_MAXISRCTDATA68 (MAXISRCTDATA[68], MAXISRCTDATA_OUT[68]);
  buf B_MAXISRCTDATA69 (MAXISRCTDATA[69], MAXISRCTDATA_OUT[69]);
  buf B_MAXISRCTDATA7 (MAXISRCTDATA[7], MAXISRCTDATA_OUT[7]);
  buf B_MAXISRCTDATA70 (MAXISRCTDATA[70], MAXISRCTDATA_OUT[70]);
  buf B_MAXISRCTDATA71 (MAXISRCTDATA[71], MAXISRCTDATA_OUT[71]);
  buf B_MAXISRCTDATA72 (MAXISRCTDATA[72], MAXISRCTDATA_OUT[72]);
  buf B_MAXISRCTDATA73 (MAXISRCTDATA[73], MAXISRCTDATA_OUT[73]);
  buf B_MAXISRCTDATA74 (MAXISRCTDATA[74], MAXISRCTDATA_OUT[74]);
  buf B_MAXISRCTDATA75 (MAXISRCTDATA[75], MAXISRCTDATA_OUT[75]);
  buf B_MAXISRCTDATA76 (MAXISRCTDATA[76], MAXISRCTDATA_OUT[76]);
  buf B_MAXISRCTDATA77 (MAXISRCTDATA[77], MAXISRCTDATA_OUT[77]);
  buf B_MAXISRCTDATA78 (MAXISRCTDATA[78], MAXISRCTDATA_OUT[78]);
  buf B_MAXISRCTDATA79 (MAXISRCTDATA[79], MAXISRCTDATA_OUT[79]);
  buf B_MAXISRCTDATA8 (MAXISRCTDATA[8], MAXISRCTDATA_OUT[8]);
  buf B_MAXISRCTDATA80 (MAXISRCTDATA[80], MAXISRCTDATA_OUT[80]);
  buf B_MAXISRCTDATA81 (MAXISRCTDATA[81], MAXISRCTDATA_OUT[81]);
  buf B_MAXISRCTDATA82 (MAXISRCTDATA[82], MAXISRCTDATA_OUT[82]);
  buf B_MAXISRCTDATA83 (MAXISRCTDATA[83], MAXISRCTDATA_OUT[83]);
  buf B_MAXISRCTDATA84 (MAXISRCTDATA[84], MAXISRCTDATA_OUT[84]);
  buf B_MAXISRCTDATA85 (MAXISRCTDATA[85], MAXISRCTDATA_OUT[85]);
  buf B_MAXISRCTDATA86 (MAXISRCTDATA[86], MAXISRCTDATA_OUT[86]);
  buf B_MAXISRCTDATA87 (MAXISRCTDATA[87], MAXISRCTDATA_OUT[87]);
  buf B_MAXISRCTDATA88 (MAXISRCTDATA[88], MAXISRCTDATA_OUT[88]);
  buf B_MAXISRCTDATA89 (MAXISRCTDATA[89], MAXISRCTDATA_OUT[89]);
  buf B_MAXISRCTDATA9 (MAXISRCTDATA[9], MAXISRCTDATA_OUT[9]);
  buf B_MAXISRCTDATA90 (MAXISRCTDATA[90], MAXISRCTDATA_OUT[90]);
  buf B_MAXISRCTDATA91 (MAXISRCTDATA[91], MAXISRCTDATA_OUT[91]);
  buf B_MAXISRCTDATA92 (MAXISRCTDATA[92], MAXISRCTDATA_OUT[92]);
  buf B_MAXISRCTDATA93 (MAXISRCTDATA[93], MAXISRCTDATA_OUT[93]);
  buf B_MAXISRCTDATA94 (MAXISRCTDATA[94], MAXISRCTDATA_OUT[94]);
  buf B_MAXISRCTDATA95 (MAXISRCTDATA[95], MAXISRCTDATA_OUT[95]);
  buf B_MAXISRCTDATA96 (MAXISRCTDATA[96], MAXISRCTDATA_OUT[96]);
  buf B_MAXISRCTDATA97 (MAXISRCTDATA[97], MAXISRCTDATA_OUT[97]);
  buf B_MAXISRCTDATA98 (MAXISRCTDATA[98], MAXISRCTDATA_OUT[98]);
  buf B_MAXISRCTDATA99 (MAXISRCTDATA[99], MAXISRCTDATA_OUT[99]);
  buf B_MAXISRCTKEEP0 (MAXISRCTKEEP[0], MAXISRCTKEEP_OUT[0]);
  buf B_MAXISRCTKEEP1 (MAXISRCTKEEP[1], MAXISRCTKEEP_OUT[1]);
  buf B_MAXISRCTKEEP2 (MAXISRCTKEEP[2], MAXISRCTKEEP_OUT[2]);
  buf B_MAXISRCTKEEP3 (MAXISRCTKEEP[3], MAXISRCTKEEP_OUT[3]);
  buf B_MAXISRCTKEEP4 (MAXISRCTKEEP[4], MAXISRCTKEEP_OUT[4]);
  buf B_MAXISRCTKEEP5 (MAXISRCTKEEP[5], MAXISRCTKEEP_OUT[5]);
  buf B_MAXISRCTKEEP6 (MAXISRCTKEEP[6], MAXISRCTKEEP_OUT[6]);
  buf B_MAXISRCTKEEP7 (MAXISRCTKEEP[7], MAXISRCTKEEP_OUT[7]);
  buf B_MAXISRCTLAST (MAXISRCTLAST, MAXISRCTLAST_OUT);
  buf B_MAXISRCTUSER0 (MAXISRCTUSER[0], MAXISRCTUSER_OUT[0]);
  buf B_MAXISRCTUSER1 (MAXISRCTUSER[1], MAXISRCTUSER_OUT[1]);
  buf B_MAXISRCTUSER10 (MAXISRCTUSER[10], MAXISRCTUSER_OUT[10]);
  buf B_MAXISRCTUSER11 (MAXISRCTUSER[11], MAXISRCTUSER_OUT[11]);
  buf B_MAXISRCTUSER12 (MAXISRCTUSER[12], MAXISRCTUSER_OUT[12]);
  buf B_MAXISRCTUSER13 (MAXISRCTUSER[13], MAXISRCTUSER_OUT[13]);
  buf B_MAXISRCTUSER14 (MAXISRCTUSER[14], MAXISRCTUSER_OUT[14]);
  buf B_MAXISRCTUSER15 (MAXISRCTUSER[15], MAXISRCTUSER_OUT[15]);
  buf B_MAXISRCTUSER16 (MAXISRCTUSER[16], MAXISRCTUSER_OUT[16]);
  buf B_MAXISRCTUSER17 (MAXISRCTUSER[17], MAXISRCTUSER_OUT[17]);
  buf B_MAXISRCTUSER18 (MAXISRCTUSER[18], MAXISRCTUSER_OUT[18]);
  buf B_MAXISRCTUSER19 (MAXISRCTUSER[19], MAXISRCTUSER_OUT[19]);
  buf B_MAXISRCTUSER2 (MAXISRCTUSER[2], MAXISRCTUSER_OUT[2]);
  buf B_MAXISRCTUSER20 (MAXISRCTUSER[20], MAXISRCTUSER_OUT[20]);
  buf B_MAXISRCTUSER21 (MAXISRCTUSER[21], MAXISRCTUSER_OUT[21]);
  buf B_MAXISRCTUSER22 (MAXISRCTUSER[22], MAXISRCTUSER_OUT[22]);
  buf B_MAXISRCTUSER23 (MAXISRCTUSER[23], MAXISRCTUSER_OUT[23]);
  buf B_MAXISRCTUSER24 (MAXISRCTUSER[24], MAXISRCTUSER_OUT[24]);
  buf B_MAXISRCTUSER25 (MAXISRCTUSER[25], MAXISRCTUSER_OUT[25]);
  buf B_MAXISRCTUSER26 (MAXISRCTUSER[26], MAXISRCTUSER_OUT[26]);
  buf B_MAXISRCTUSER27 (MAXISRCTUSER[27], MAXISRCTUSER_OUT[27]);
  buf B_MAXISRCTUSER28 (MAXISRCTUSER[28], MAXISRCTUSER_OUT[28]);
  buf B_MAXISRCTUSER29 (MAXISRCTUSER[29], MAXISRCTUSER_OUT[29]);
  buf B_MAXISRCTUSER3 (MAXISRCTUSER[3], MAXISRCTUSER_OUT[3]);
  buf B_MAXISRCTUSER30 (MAXISRCTUSER[30], MAXISRCTUSER_OUT[30]);
  buf B_MAXISRCTUSER31 (MAXISRCTUSER[31], MAXISRCTUSER_OUT[31]);
  buf B_MAXISRCTUSER32 (MAXISRCTUSER[32], MAXISRCTUSER_OUT[32]);
  buf B_MAXISRCTUSER33 (MAXISRCTUSER[33], MAXISRCTUSER_OUT[33]);
  buf B_MAXISRCTUSER34 (MAXISRCTUSER[34], MAXISRCTUSER_OUT[34]);
  buf B_MAXISRCTUSER35 (MAXISRCTUSER[35], MAXISRCTUSER_OUT[35]);
  buf B_MAXISRCTUSER36 (MAXISRCTUSER[36], MAXISRCTUSER_OUT[36]);
  buf B_MAXISRCTUSER37 (MAXISRCTUSER[37], MAXISRCTUSER_OUT[37]);
  buf B_MAXISRCTUSER38 (MAXISRCTUSER[38], MAXISRCTUSER_OUT[38]);
  buf B_MAXISRCTUSER39 (MAXISRCTUSER[39], MAXISRCTUSER_OUT[39]);
  buf B_MAXISRCTUSER4 (MAXISRCTUSER[4], MAXISRCTUSER_OUT[4]);
  buf B_MAXISRCTUSER40 (MAXISRCTUSER[40], MAXISRCTUSER_OUT[40]);
  buf B_MAXISRCTUSER41 (MAXISRCTUSER[41], MAXISRCTUSER_OUT[41]);
  buf B_MAXISRCTUSER42 (MAXISRCTUSER[42], MAXISRCTUSER_OUT[42]);
  buf B_MAXISRCTUSER43 (MAXISRCTUSER[43], MAXISRCTUSER_OUT[43]);
  buf B_MAXISRCTUSER44 (MAXISRCTUSER[44], MAXISRCTUSER_OUT[44]);
  buf B_MAXISRCTUSER45 (MAXISRCTUSER[45], MAXISRCTUSER_OUT[45]);
  buf B_MAXISRCTUSER46 (MAXISRCTUSER[46], MAXISRCTUSER_OUT[46]);
  buf B_MAXISRCTUSER47 (MAXISRCTUSER[47], MAXISRCTUSER_OUT[47]);
  buf B_MAXISRCTUSER48 (MAXISRCTUSER[48], MAXISRCTUSER_OUT[48]);
  buf B_MAXISRCTUSER49 (MAXISRCTUSER[49], MAXISRCTUSER_OUT[49]);
  buf B_MAXISRCTUSER5 (MAXISRCTUSER[5], MAXISRCTUSER_OUT[5]);
  buf B_MAXISRCTUSER50 (MAXISRCTUSER[50], MAXISRCTUSER_OUT[50]);
  buf B_MAXISRCTUSER51 (MAXISRCTUSER[51], MAXISRCTUSER_OUT[51]);
  buf B_MAXISRCTUSER52 (MAXISRCTUSER[52], MAXISRCTUSER_OUT[52]);
  buf B_MAXISRCTUSER53 (MAXISRCTUSER[53], MAXISRCTUSER_OUT[53]);
  buf B_MAXISRCTUSER54 (MAXISRCTUSER[54], MAXISRCTUSER_OUT[54]);
  buf B_MAXISRCTUSER55 (MAXISRCTUSER[55], MAXISRCTUSER_OUT[55]);
  buf B_MAXISRCTUSER56 (MAXISRCTUSER[56], MAXISRCTUSER_OUT[56]);
  buf B_MAXISRCTUSER57 (MAXISRCTUSER[57], MAXISRCTUSER_OUT[57]);
  buf B_MAXISRCTUSER58 (MAXISRCTUSER[58], MAXISRCTUSER_OUT[58]);
  buf B_MAXISRCTUSER59 (MAXISRCTUSER[59], MAXISRCTUSER_OUT[59]);
  buf B_MAXISRCTUSER6 (MAXISRCTUSER[6], MAXISRCTUSER_OUT[6]);
  buf B_MAXISRCTUSER60 (MAXISRCTUSER[60], MAXISRCTUSER_OUT[60]);
  buf B_MAXISRCTUSER61 (MAXISRCTUSER[61], MAXISRCTUSER_OUT[61]);
  buf B_MAXISRCTUSER62 (MAXISRCTUSER[62], MAXISRCTUSER_OUT[62]);
  buf B_MAXISRCTUSER63 (MAXISRCTUSER[63], MAXISRCTUSER_OUT[63]);
  buf B_MAXISRCTUSER64 (MAXISRCTUSER[64], MAXISRCTUSER_OUT[64]);
  buf B_MAXISRCTUSER65 (MAXISRCTUSER[65], MAXISRCTUSER_OUT[65]);
  buf B_MAXISRCTUSER66 (MAXISRCTUSER[66], MAXISRCTUSER_OUT[66]);
  buf B_MAXISRCTUSER67 (MAXISRCTUSER[67], MAXISRCTUSER_OUT[67]);
  buf B_MAXISRCTUSER68 (MAXISRCTUSER[68], MAXISRCTUSER_OUT[68]);
  buf B_MAXISRCTUSER69 (MAXISRCTUSER[69], MAXISRCTUSER_OUT[69]);
  buf B_MAXISRCTUSER7 (MAXISRCTUSER[7], MAXISRCTUSER_OUT[7]);
  buf B_MAXISRCTUSER70 (MAXISRCTUSER[70], MAXISRCTUSER_OUT[70]);
  buf B_MAXISRCTUSER71 (MAXISRCTUSER[71], MAXISRCTUSER_OUT[71]);
  buf B_MAXISRCTUSER72 (MAXISRCTUSER[72], MAXISRCTUSER_OUT[72]);
  buf B_MAXISRCTUSER73 (MAXISRCTUSER[73], MAXISRCTUSER_OUT[73]);
  buf B_MAXISRCTUSER74 (MAXISRCTUSER[74], MAXISRCTUSER_OUT[74]);
  buf B_MAXISRCTUSER8 (MAXISRCTUSER[8], MAXISRCTUSER_OUT[8]);
  buf B_MAXISRCTUSER9 (MAXISRCTUSER[9], MAXISRCTUSER_OUT[9]);
  buf B_MAXISRCTVALID (MAXISRCTVALID, MAXISRCTVALID_OUT);
  buf B_MICOMPLETIONRAMREADADDRESSAL0 (MICOMPLETIONRAMREADADDRESSAL[0], MICOMPLETIONRAMREADADDRESSAL_OUT[0]);
  buf B_MICOMPLETIONRAMREADADDRESSAL1 (MICOMPLETIONRAMREADADDRESSAL[1], MICOMPLETIONRAMREADADDRESSAL_OUT[1]);
  buf B_MICOMPLETIONRAMREADADDRESSAL2 (MICOMPLETIONRAMREADADDRESSAL[2], MICOMPLETIONRAMREADADDRESSAL_OUT[2]);
  buf B_MICOMPLETIONRAMREADADDRESSAL3 (MICOMPLETIONRAMREADADDRESSAL[3], MICOMPLETIONRAMREADADDRESSAL_OUT[3]);
  buf B_MICOMPLETIONRAMREADADDRESSAL4 (MICOMPLETIONRAMREADADDRESSAL[4], MICOMPLETIONRAMREADADDRESSAL_OUT[4]);
  buf B_MICOMPLETIONRAMREADADDRESSAL5 (MICOMPLETIONRAMREADADDRESSAL[5], MICOMPLETIONRAMREADADDRESSAL_OUT[5]);
  buf B_MICOMPLETIONRAMREADADDRESSAL6 (MICOMPLETIONRAMREADADDRESSAL[6], MICOMPLETIONRAMREADADDRESSAL_OUT[6]);
  buf B_MICOMPLETIONRAMREADADDRESSAL7 (MICOMPLETIONRAMREADADDRESSAL[7], MICOMPLETIONRAMREADADDRESSAL_OUT[7]);
  buf B_MICOMPLETIONRAMREADADDRESSAL8 (MICOMPLETIONRAMREADADDRESSAL[8], MICOMPLETIONRAMREADADDRESSAL_OUT[8]);
  buf B_MICOMPLETIONRAMREADADDRESSAL9 (MICOMPLETIONRAMREADADDRESSAL[9], MICOMPLETIONRAMREADADDRESSAL_OUT[9]);
  buf B_MICOMPLETIONRAMREADADDRESSAU0 (MICOMPLETIONRAMREADADDRESSAU[0], MICOMPLETIONRAMREADADDRESSAU_OUT[0]);
  buf B_MICOMPLETIONRAMREADADDRESSAU1 (MICOMPLETIONRAMREADADDRESSAU[1], MICOMPLETIONRAMREADADDRESSAU_OUT[1]);
  buf B_MICOMPLETIONRAMREADADDRESSAU2 (MICOMPLETIONRAMREADADDRESSAU[2], MICOMPLETIONRAMREADADDRESSAU_OUT[2]);
  buf B_MICOMPLETIONRAMREADADDRESSAU3 (MICOMPLETIONRAMREADADDRESSAU[3], MICOMPLETIONRAMREADADDRESSAU_OUT[3]);
  buf B_MICOMPLETIONRAMREADADDRESSAU4 (MICOMPLETIONRAMREADADDRESSAU[4], MICOMPLETIONRAMREADADDRESSAU_OUT[4]);
  buf B_MICOMPLETIONRAMREADADDRESSAU5 (MICOMPLETIONRAMREADADDRESSAU[5], MICOMPLETIONRAMREADADDRESSAU_OUT[5]);
  buf B_MICOMPLETIONRAMREADADDRESSAU6 (MICOMPLETIONRAMREADADDRESSAU[6], MICOMPLETIONRAMREADADDRESSAU_OUT[6]);
  buf B_MICOMPLETIONRAMREADADDRESSAU7 (MICOMPLETIONRAMREADADDRESSAU[7], MICOMPLETIONRAMREADADDRESSAU_OUT[7]);
  buf B_MICOMPLETIONRAMREADADDRESSAU8 (MICOMPLETIONRAMREADADDRESSAU[8], MICOMPLETIONRAMREADADDRESSAU_OUT[8]);
  buf B_MICOMPLETIONRAMREADADDRESSAU9 (MICOMPLETIONRAMREADADDRESSAU[9], MICOMPLETIONRAMREADADDRESSAU_OUT[9]);
  buf B_MICOMPLETIONRAMREADADDRESSBL0 (MICOMPLETIONRAMREADADDRESSBL[0], MICOMPLETIONRAMREADADDRESSBL_OUT[0]);
  buf B_MICOMPLETIONRAMREADADDRESSBL1 (MICOMPLETIONRAMREADADDRESSBL[1], MICOMPLETIONRAMREADADDRESSBL_OUT[1]);
  buf B_MICOMPLETIONRAMREADADDRESSBL2 (MICOMPLETIONRAMREADADDRESSBL[2], MICOMPLETIONRAMREADADDRESSBL_OUT[2]);
  buf B_MICOMPLETIONRAMREADADDRESSBL3 (MICOMPLETIONRAMREADADDRESSBL[3], MICOMPLETIONRAMREADADDRESSBL_OUT[3]);
  buf B_MICOMPLETIONRAMREADADDRESSBL4 (MICOMPLETIONRAMREADADDRESSBL[4], MICOMPLETIONRAMREADADDRESSBL_OUT[4]);
  buf B_MICOMPLETIONRAMREADADDRESSBL5 (MICOMPLETIONRAMREADADDRESSBL[5], MICOMPLETIONRAMREADADDRESSBL_OUT[5]);
  buf B_MICOMPLETIONRAMREADADDRESSBL6 (MICOMPLETIONRAMREADADDRESSBL[6], MICOMPLETIONRAMREADADDRESSBL_OUT[6]);
  buf B_MICOMPLETIONRAMREADADDRESSBL7 (MICOMPLETIONRAMREADADDRESSBL[7], MICOMPLETIONRAMREADADDRESSBL_OUT[7]);
  buf B_MICOMPLETIONRAMREADADDRESSBL8 (MICOMPLETIONRAMREADADDRESSBL[8], MICOMPLETIONRAMREADADDRESSBL_OUT[8]);
  buf B_MICOMPLETIONRAMREADADDRESSBL9 (MICOMPLETIONRAMREADADDRESSBL[9], MICOMPLETIONRAMREADADDRESSBL_OUT[9]);
  buf B_MICOMPLETIONRAMREADADDRESSBU0 (MICOMPLETIONRAMREADADDRESSBU[0], MICOMPLETIONRAMREADADDRESSBU_OUT[0]);
  buf B_MICOMPLETIONRAMREADADDRESSBU1 (MICOMPLETIONRAMREADADDRESSBU[1], MICOMPLETIONRAMREADADDRESSBU_OUT[1]);
  buf B_MICOMPLETIONRAMREADADDRESSBU2 (MICOMPLETIONRAMREADADDRESSBU[2], MICOMPLETIONRAMREADADDRESSBU_OUT[2]);
  buf B_MICOMPLETIONRAMREADADDRESSBU3 (MICOMPLETIONRAMREADADDRESSBU[3], MICOMPLETIONRAMREADADDRESSBU_OUT[3]);
  buf B_MICOMPLETIONRAMREADADDRESSBU4 (MICOMPLETIONRAMREADADDRESSBU[4], MICOMPLETIONRAMREADADDRESSBU_OUT[4]);
  buf B_MICOMPLETIONRAMREADADDRESSBU5 (MICOMPLETIONRAMREADADDRESSBU[5], MICOMPLETIONRAMREADADDRESSBU_OUT[5]);
  buf B_MICOMPLETIONRAMREADADDRESSBU6 (MICOMPLETIONRAMREADADDRESSBU[6], MICOMPLETIONRAMREADADDRESSBU_OUT[6]);
  buf B_MICOMPLETIONRAMREADADDRESSBU7 (MICOMPLETIONRAMREADADDRESSBU[7], MICOMPLETIONRAMREADADDRESSBU_OUT[7]);
  buf B_MICOMPLETIONRAMREADADDRESSBU8 (MICOMPLETIONRAMREADADDRESSBU[8], MICOMPLETIONRAMREADADDRESSBU_OUT[8]);
  buf B_MICOMPLETIONRAMREADADDRESSBU9 (MICOMPLETIONRAMREADADDRESSBU[9], MICOMPLETIONRAMREADADDRESSBU_OUT[9]);
  buf B_MICOMPLETIONRAMREADENABLEL0 (MICOMPLETIONRAMREADENABLEL[0], MICOMPLETIONRAMREADENABLEL_OUT[0]);
  buf B_MICOMPLETIONRAMREADENABLEL1 (MICOMPLETIONRAMREADENABLEL[1], MICOMPLETIONRAMREADENABLEL_OUT[1]);
  buf B_MICOMPLETIONRAMREADENABLEL2 (MICOMPLETIONRAMREADENABLEL[2], MICOMPLETIONRAMREADENABLEL_OUT[2]);
  buf B_MICOMPLETIONRAMREADENABLEL3 (MICOMPLETIONRAMREADENABLEL[3], MICOMPLETIONRAMREADENABLEL_OUT[3]);
  buf B_MICOMPLETIONRAMREADENABLEU0 (MICOMPLETIONRAMREADENABLEU[0], MICOMPLETIONRAMREADENABLEU_OUT[0]);
  buf B_MICOMPLETIONRAMREADENABLEU1 (MICOMPLETIONRAMREADENABLEU[1], MICOMPLETIONRAMREADENABLEU_OUT[1]);
  buf B_MICOMPLETIONRAMREADENABLEU2 (MICOMPLETIONRAMREADENABLEU[2], MICOMPLETIONRAMREADENABLEU_OUT[2]);
  buf B_MICOMPLETIONRAMREADENABLEU3 (MICOMPLETIONRAMREADENABLEU[3], MICOMPLETIONRAMREADENABLEU_OUT[3]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAL0 (MICOMPLETIONRAMWRITEADDRESSAL[0], MICOMPLETIONRAMWRITEADDRESSAL_OUT[0]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAL1 (MICOMPLETIONRAMWRITEADDRESSAL[1], MICOMPLETIONRAMWRITEADDRESSAL_OUT[1]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAL2 (MICOMPLETIONRAMWRITEADDRESSAL[2], MICOMPLETIONRAMWRITEADDRESSAL_OUT[2]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAL3 (MICOMPLETIONRAMWRITEADDRESSAL[3], MICOMPLETIONRAMWRITEADDRESSAL_OUT[3]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAL4 (MICOMPLETIONRAMWRITEADDRESSAL[4], MICOMPLETIONRAMWRITEADDRESSAL_OUT[4]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAL5 (MICOMPLETIONRAMWRITEADDRESSAL[5], MICOMPLETIONRAMWRITEADDRESSAL_OUT[5]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAL6 (MICOMPLETIONRAMWRITEADDRESSAL[6], MICOMPLETIONRAMWRITEADDRESSAL_OUT[6]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAL7 (MICOMPLETIONRAMWRITEADDRESSAL[7], MICOMPLETIONRAMWRITEADDRESSAL_OUT[7]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAL8 (MICOMPLETIONRAMWRITEADDRESSAL[8], MICOMPLETIONRAMWRITEADDRESSAL_OUT[8]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAL9 (MICOMPLETIONRAMWRITEADDRESSAL[9], MICOMPLETIONRAMWRITEADDRESSAL_OUT[9]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAU0 (MICOMPLETIONRAMWRITEADDRESSAU[0], MICOMPLETIONRAMWRITEADDRESSAU_OUT[0]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAU1 (MICOMPLETIONRAMWRITEADDRESSAU[1], MICOMPLETIONRAMWRITEADDRESSAU_OUT[1]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAU2 (MICOMPLETIONRAMWRITEADDRESSAU[2], MICOMPLETIONRAMWRITEADDRESSAU_OUT[2]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAU3 (MICOMPLETIONRAMWRITEADDRESSAU[3], MICOMPLETIONRAMWRITEADDRESSAU_OUT[3]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAU4 (MICOMPLETIONRAMWRITEADDRESSAU[4], MICOMPLETIONRAMWRITEADDRESSAU_OUT[4]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAU5 (MICOMPLETIONRAMWRITEADDRESSAU[5], MICOMPLETIONRAMWRITEADDRESSAU_OUT[5]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAU6 (MICOMPLETIONRAMWRITEADDRESSAU[6], MICOMPLETIONRAMWRITEADDRESSAU_OUT[6]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAU7 (MICOMPLETIONRAMWRITEADDRESSAU[7], MICOMPLETIONRAMWRITEADDRESSAU_OUT[7]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAU8 (MICOMPLETIONRAMWRITEADDRESSAU[8], MICOMPLETIONRAMWRITEADDRESSAU_OUT[8]);
  buf B_MICOMPLETIONRAMWRITEADDRESSAU9 (MICOMPLETIONRAMWRITEADDRESSAU[9], MICOMPLETIONRAMWRITEADDRESSAU_OUT[9]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBL0 (MICOMPLETIONRAMWRITEADDRESSBL[0], MICOMPLETIONRAMWRITEADDRESSBL_OUT[0]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBL1 (MICOMPLETIONRAMWRITEADDRESSBL[1], MICOMPLETIONRAMWRITEADDRESSBL_OUT[1]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBL2 (MICOMPLETIONRAMWRITEADDRESSBL[2], MICOMPLETIONRAMWRITEADDRESSBL_OUT[2]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBL3 (MICOMPLETIONRAMWRITEADDRESSBL[3], MICOMPLETIONRAMWRITEADDRESSBL_OUT[3]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBL4 (MICOMPLETIONRAMWRITEADDRESSBL[4], MICOMPLETIONRAMWRITEADDRESSBL_OUT[4]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBL5 (MICOMPLETIONRAMWRITEADDRESSBL[5], MICOMPLETIONRAMWRITEADDRESSBL_OUT[5]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBL6 (MICOMPLETIONRAMWRITEADDRESSBL[6], MICOMPLETIONRAMWRITEADDRESSBL_OUT[6]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBL7 (MICOMPLETIONRAMWRITEADDRESSBL[7], MICOMPLETIONRAMWRITEADDRESSBL_OUT[7]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBL8 (MICOMPLETIONRAMWRITEADDRESSBL[8], MICOMPLETIONRAMWRITEADDRESSBL_OUT[8]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBL9 (MICOMPLETIONRAMWRITEADDRESSBL[9], MICOMPLETIONRAMWRITEADDRESSBL_OUT[9]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBU0 (MICOMPLETIONRAMWRITEADDRESSBU[0], MICOMPLETIONRAMWRITEADDRESSBU_OUT[0]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBU1 (MICOMPLETIONRAMWRITEADDRESSBU[1], MICOMPLETIONRAMWRITEADDRESSBU_OUT[1]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBU2 (MICOMPLETIONRAMWRITEADDRESSBU[2], MICOMPLETIONRAMWRITEADDRESSBU_OUT[2]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBU3 (MICOMPLETIONRAMWRITEADDRESSBU[3], MICOMPLETIONRAMWRITEADDRESSBU_OUT[3]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBU4 (MICOMPLETIONRAMWRITEADDRESSBU[4], MICOMPLETIONRAMWRITEADDRESSBU_OUT[4]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBU5 (MICOMPLETIONRAMWRITEADDRESSBU[5], MICOMPLETIONRAMWRITEADDRESSBU_OUT[5]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBU6 (MICOMPLETIONRAMWRITEADDRESSBU[6], MICOMPLETIONRAMWRITEADDRESSBU_OUT[6]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBU7 (MICOMPLETIONRAMWRITEADDRESSBU[7], MICOMPLETIONRAMWRITEADDRESSBU_OUT[7]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBU8 (MICOMPLETIONRAMWRITEADDRESSBU[8], MICOMPLETIONRAMWRITEADDRESSBU_OUT[8]);
  buf B_MICOMPLETIONRAMWRITEADDRESSBU9 (MICOMPLETIONRAMWRITEADDRESSBU[9], MICOMPLETIONRAMWRITEADDRESSBU_OUT[9]);
  buf B_MICOMPLETIONRAMWRITEDATAL0 (MICOMPLETIONRAMWRITEDATAL[0], MICOMPLETIONRAMWRITEDATAL_OUT[0]);
  buf B_MICOMPLETIONRAMWRITEDATAL1 (MICOMPLETIONRAMWRITEDATAL[1], MICOMPLETIONRAMWRITEDATAL_OUT[1]);
  buf B_MICOMPLETIONRAMWRITEDATAL10 (MICOMPLETIONRAMWRITEDATAL[10], MICOMPLETIONRAMWRITEDATAL_OUT[10]);
  buf B_MICOMPLETIONRAMWRITEDATAL11 (MICOMPLETIONRAMWRITEDATAL[11], MICOMPLETIONRAMWRITEDATAL_OUT[11]);
  buf B_MICOMPLETIONRAMWRITEDATAL12 (MICOMPLETIONRAMWRITEDATAL[12], MICOMPLETIONRAMWRITEDATAL_OUT[12]);
  buf B_MICOMPLETIONRAMWRITEDATAL13 (MICOMPLETIONRAMWRITEDATAL[13], MICOMPLETIONRAMWRITEDATAL_OUT[13]);
  buf B_MICOMPLETIONRAMWRITEDATAL14 (MICOMPLETIONRAMWRITEDATAL[14], MICOMPLETIONRAMWRITEDATAL_OUT[14]);
  buf B_MICOMPLETIONRAMWRITEDATAL15 (MICOMPLETIONRAMWRITEDATAL[15], MICOMPLETIONRAMWRITEDATAL_OUT[15]);
  buf B_MICOMPLETIONRAMWRITEDATAL16 (MICOMPLETIONRAMWRITEDATAL[16], MICOMPLETIONRAMWRITEDATAL_OUT[16]);
  buf B_MICOMPLETIONRAMWRITEDATAL17 (MICOMPLETIONRAMWRITEDATAL[17], MICOMPLETIONRAMWRITEDATAL_OUT[17]);
  buf B_MICOMPLETIONRAMWRITEDATAL18 (MICOMPLETIONRAMWRITEDATAL[18], MICOMPLETIONRAMWRITEDATAL_OUT[18]);
  buf B_MICOMPLETIONRAMWRITEDATAL19 (MICOMPLETIONRAMWRITEDATAL[19], MICOMPLETIONRAMWRITEDATAL_OUT[19]);
  buf B_MICOMPLETIONRAMWRITEDATAL2 (MICOMPLETIONRAMWRITEDATAL[2], MICOMPLETIONRAMWRITEDATAL_OUT[2]);
  buf B_MICOMPLETIONRAMWRITEDATAL20 (MICOMPLETIONRAMWRITEDATAL[20], MICOMPLETIONRAMWRITEDATAL_OUT[20]);
  buf B_MICOMPLETIONRAMWRITEDATAL21 (MICOMPLETIONRAMWRITEDATAL[21], MICOMPLETIONRAMWRITEDATAL_OUT[21]);
  buf B_MICOMPLETIONRAMWRITEDATAL22 (MICOMPLETIONRAMWRITEDATAL[22], MICOMPLETIONRAMWRITEDATAL_OUT[22]);
  buf B_MICOMPLETIONRAMWRITEDATAL23 (MICOMPLETIONRAMWRITEDATAL[23], MICOMPLETIONRAMWRITEDATAL_OUT[23]);
  buf B_MICOMPLETIONRAMWRITEDATAL24 (MICOMPLETIONRAMWRITEDATAL[24], MICOMPLETIONRAMWRITEDATAL_OUT[24]);
  buf B_MICOMPLETIONRAMWRITEDATAL25 (MICOMPLETIONRAMWRITEDATAL[25], MICOMPLETIONRAMWRITEDATAL_OUT[25]);
  buf B_MICOMPLETIONRAMWRITEDATAL26 (MICOMPLETIONRAMWRITEDATAL[26], MICOMPLETIONRAMWRITEDATAL_OUT[26]);
  buf B_MICOMPLETIONRAMWRITEDATAL27 (MICOMPLETIONRAMWRITEDATAL[27], MICOMPLETIONRAMWRITEDATAL_OUT[27]);
  buf B_MICOMPLETIONRAMWRITEDATAL28 (MICOMPLETIONRAMWRITEDATAL[28], MICOMPLETIONRAMWRITEDATAL_OUT[28]);
  buf B_MICOMPLETIONRAMWRITEDATAL29 (MICOMPLETIONRAMWRITEDATAL[29], MICOMPLETIONRAMWRITEDATAL_OUT[29]);
  buf B_MICOMPLETIONRAMWRITEDATAL3 (MICOMPLETIONRAMWRITEDATAL[3], MICOMPLETIONRAMWRITEDATAL_OUT[3]);
  buf B_MICOMPLETIONRAMWRITEDATAL30 (MICOMPLETIONRAMWRITEDATAL[30], MICOMPLETIONRAMWRITEDATAL_OUT[30]);
  buf B_MICOMPLETIONRAMWRITEDATAL31 (MICOMPLETIONRAMWRITEDATAL[31], MICOMPLETIONRAMWRITEDATAL_OUT[31]);
  buf B_MICOMPLETIONRAMWRITEDATAL32 (MICOMPLETIONRAMWRITEDATAL[32], MICOMPLETIONRAMWRITEDATAL_OUT[32]);
  buf B_MICOMPLETIONRAMWRITEDATAL33 (MICOMPLETIONRAMWRITEDATAL[33], MICOMPLETIONRAMWRITEDATAL_OUT[33]);
  buf B_MICOMPLETIONRAMWRITEDATAL34 (MICOMPLETIONRAMWRITEDATAL[34], MICOMPLETIONRAMWRITEDATAL_OUT[34]);
  buf B_MICOMPLETIONRAMWRITEDATAL35 (MICOMPLETIONRAMWRITEDATAL[35], MICOMPLETIONRAMWRITEDATAL_OUT[35]);
  buf B_MICOMPLETIONRAMWRITEDATAL36 (MICOMPLETIONRAMWRITEDATAL[36], MICOMPLETIONRAMWRITEDATAL_OUT[36]);
  buf B_MICOMPLETIONRAMWRITEDATAL37 (MICOMPLETIONRAMWRITEDATAL[37], MICOMPLETIONRAMWRITEDATAL_OUT[37]);
  buf B_MICOMPLETIONRAMWRITEDATAL38 (MICOMPLETIONRAMWRITEDATAL[38], MICOMPLETIONRAMWRITEDATAL_OUT[38]);
  buf B_MICOMPLETIONRAMWRITEDATAL39 (MICOMPLETIONRAMWRITEDATAL[39], MICOMPLETIONRAMWRITEDATAL_OUT[39]);
  buf B_MICOMPLETIONRAMWRITEDATAL4 (MICOMPLETIONRAMWRITEDATAL[4], MICOMPLETIONRAMWRITEDATAL_OUT[4]);
  buf B_MICOMPLETIONRAMWRITEDATAL40 (MICOMPLETIONRAMWRITEDATAL[40], MICOMPLETIONRAMWRITEDATAL_OUT[40]);
  buf B_MICOMPLETIONRAMWRITEDATAL41 (MICOMPLETIONRAMWRITEDATAL[41], MICOMPLETIONRAMWRITEDATAL_OUT[41]);
  buf B_MICOMPLETIONRAMWRITEDATAL42 (MICOMPLETIONRAMWRITEDATAL[42], MICOMPLETIONRAMWRITEDATAL_OUT[42]);
  buf B_MICOMPLETIONRAMWRITEDATAL43 (MICOMPLETIONRAMWRITEDATAL[43], MICOMPLETIONRAMWRITEDATAL_OUT[43]);
  buf B_MICOMPLETIONRAMWRITEDATAL44 (MICOMPLETIONRAMWRITEDATAL[44], MICOMPLETIONRAMWRITEDATAL_OUT[44]);
  buf B_MICOMPLETIONRAMWRITEDATAL45 (MICOMPLETIONRAMWRITEDATAL[45], MICOMPLETIONRAMWRITEDATAL_OUT[45]);
  buf B_MICOMPLETIONRAMWRITEDATAL46 (MICOMPLETIONRAMWRITEDATAL[46], MICOMPLETIONRAMWRITEDATAL_OUT[46]);
  buf B_MICOMPLETIONRAMWRITEDATAL47 (MICOMPLETIONRAMWRITEDATAL[47], MICOMPLETIONRAMWRITEDATAL_OUT[47]);
  buf B_MICOMPLETIONRAMWRITEDATAL48 (MICOMPLETIONRAMWRITEDATAL[48], MICOMPLETIONRAMWRITEDATAL_OUT[48]);
  buf B_MICOMPLETIONRAMWRITEDATAL49 (MICOMPLETIONRAMWRITEDATAL[49], MICOMPLETIONRAMWRITEDATAL_OUT[49]);
  buf B_MICOMPLETIONRAMWRITEDATAL5 (MICOMPLETIONRAMWRITEDATAL[5], MICOMPLETIONRAMWRITEDATAL_OUT[5]);
  buf B_MICOMPLETIONRAMWRITEDATAL50 (MICOMPLETIONRAMWRITEDATAL[50], MICOMPLETIONRAMWRITEDATAL_OUT[50]);
  buf B_MICOMPLETIONRAMWRITEDATAL51 (MICOMPLETIONRAMWRITEDATAL[51], MICOMPLETIONRAMWRITEDATAL_OUT[51]);
  buf B_MICOMPLETIONRAMWRITEDATAL52 (MICOMPLETIONRAMWRITEDATAL[52], MICOMPLETIONRAMWRITEDATAL_OUT[52]);
  buf B_MICOMPLETIONRAMWRITEDATAL53 (MICOMPLETIONRAMWRITEDATAL[53], MICOMPLETIONRAMWRITEDATAL_OUT[53]);
  buf B_MICOMPLETIONRAMWRITEDATAL54 (MICOMPLETIONRAMWRITEDATAL[54], MICOMPLETIONRAMWRITEDATAL_OUT[54]);
  buf B_MICOMPLETIONRAMWRITEDATAL55 (MICOMPLETIONRAMWRITEDATAL[55], MICOMPLETIONRAMWRITEDATAL_OUT[55]);
  buf B_MICOMPLETIONRAMWRITEDATAL56 (MICOMPLETIONRAMWRITEDATAL[56], MICOMPLETIONRAMWRITEDATAL_OUT[56]);
  buf B_MICOMPLETIONRAMWRITEDATAL57 (MICOMPLETIONRAMWRITEDATAL[57], MICOMPLETIONRAMWRITEDATAL_OUT[57]);
  buf B_MICOMPLETIONRAMWRITEDATAL58 (MICOMPLETIONRAMWRITEDATAL[58], MICOMPLETIONRAMWRITEDATAL_OUT[58]);
  buf B_MICOMPLETIONRAMWRITEDATAL59 (MICOMPLETIONRAMWRITEDATAL[59], MICOMPLETIONRAMWRITEDATAL_OUT[59]);
  buf B_MICOMPLETIONRAMWRITEDATAL6 (MICOMPLETIONRAMWRITEDATAL[6], MICOMPLETIONRAMWRITEDATAL_OUT[6]);
  buf B_MICOMPLETIONRAMWRITEDATAL60 (MICOMPLETIONRAMWRITEDATAL[60], MICOMPLETIONRAMWRITEDATAL_OUT[60]);
  buf B_MICOMPLETIONRAMWRITEDATAL61 (MICOMPLETIONRAMWRITEDATAL[61], MICOMPLETIONRAMWRITEDATAL_OUT[61]);
  buf B_MICOMPLETIONRAMWRITEDATAL62 (MICOMPLETIONRAMWRITEDATAL[62], MICOMPLETIONRAMWRITEDATAL_OUT[62]);
  buf B_MICOMPLETIONRAMWRITEDATAL63 (MICOMPLETIONRAMWRITEDATAL[63], MICOMPLETIONRAMWRITEDATAL_OUT[63]);
  buf B_MICOMPLETIONRAMWRITEDATAL64 (MICOMPLETIONRAMWRITEDATAL[64], MICOMPLETIONRAMWRITEDATAL_OUT[64]);
  buf B_MICOMPLETIONRAMWRITEDATAL65 (MICOMPLETIONRAMWRITEDATAL[65], MICOMPLETIONRAMWRITEDATAL_OUT[65]);
  buf B_MICOMPLETIONRAMWRITEDATAL66 (MICOMPLETIONRAMWRITEDATAL[66], MICOMPLETIONRAMWRITEDATAL_OUT[66]);
  buf B_MICOMPLETIONRAMWRITEDATAL67 (MICOMPLETIONRAMWRITEDATAL[67], MICOMPLETIONRAMWRITEDATAL_OUT[67]);
  buf B_MICOMPLETIONRAMWRITEDATAL68 (MICOMPLETIONRAMWRITEDATAL[68], MICOMPLETIONRAMWRITEDATAL_OUT[68]);
  buf B_MICOMPLETIONRAMWRITEDATAL69 (MICOMPLETIONRAMWRITEDATAL[69], MICOMPLETIONRAMWRITEDATAL_OUT[69]);
  buf B_MICOMPLETIONRAMWRITEDATAL7 (MICOMPLETIONRAMWRITEDATAL[7], MICOMPLETIONRAMWRITEDATAL_OUT[7]);
  buf B_MICOMPLETIONRAMWRITEDATAL70 (MICOMPLETIONRAMWRITEDATAL[70], MICOMPLETIONRAMWRITEDATAL_OUT[70]);
  buf B_MICOMPLETIONRAMWRITEDATAL71 (MICOMPLETIONRAMWRITEDATAL[71], MICOMPLETIONRAMWRITEDATAL_OUT[71]);
  buf B_MICOMPLETIONRAMWRITEDATAL8 (MICOMPLETIONRAMWRITEDATAL[8], MICOMPLETIONRAMWRITEDATAL_OUT[8]);
  buf B_MICOMPLETIONRAMWRITEDATAL9 (MICOMPLETIONRAMWRITEDATAL[9], MICOMPLETIONRAMWRITEDATAL_OUT[9]);
  buf B_MICOMPLETIONRAMWRITEDATAU0 (MICOMPLETIONRAMWRITEDATAU[0], MICOMPLETIONRAMWRITEDATAU_OUT[0]);
  buf B_MICOMPLETIONRAMWRITEDATAU1 (MICOMPLETIONRAMWRITEDATAU[1], MICOMPLETIONRAMWRITEDATAU_OUT[1]);
  buf B_MICOMPLETIONRAMWRITEDATAU10 (MICOMPLETIONRAMWRITEDATAU[10], MICOMPLETIONRAMWRITEDATAU_OUT[10]);
  buf B_MICOMPLETIONRAMWRITEDATAU11 (MICOMPLETIONRAMWRITEDATAU[11], MICOMPLETIONRAMWRITEDATAU_OUT[11]);
  buf B_MICOMPLETIONRAMWRITEDATAU12 (MICOMPLETIONRAMWRITEDATAU[12], MICOMPLETIONRAMWRITEDATAU_OUT[12]);
  buf B_MICOMPLETIONRAMWRITEDATAU13 (MICOMPLETIONRAMWRITEDATAU[13], MICOMPLETIONRAMWRITEDATAU_OUT[13]);
  buf B_MICOMPLETIONRAMWRITEDATAU14 (MICOMPLETIONRAMWRITEDATAU[14], MICOMPLETIONRAMWRITEDATAU_OUT[14]);
  buf B_MICOMPLETIONRAMWRITEDATAU15 (MICOMPLETIONRAMWRITEDATAU[15], MICOMPLETIONRAMWRITEDATAU_OUT[15]);
  buf B_MICOMPLETIONRAMWRITEDATAU16 (MICOMPLETIONRAMWRITEDATAU[16], MICOMPLETIONRAMWRITEDATAU_OUT[16]);
  buf B_MICOMPLETIONRAMWRITEDATAU17 (MICOMPLETIONRAMWRITEDATAU[17], MICOMPLETIONRAMWRITEDATAU_OUT[17]);
  buf B_MICOMPLETIONRAMWRITEDATAU18 (MICOMPLETIONRAMWRITEDATAU[18], MICOMPLETIONRAMWRITEDATAU_OUT[18]);
  buf B_MICOMPLETIONRAMWRITEDATAU19 (MICOMPLETIONRAMWRITEDATAU[19], MICOMPLETIONRAMWRITEDATAU_OUT[19]);
  buf B_MICOMPLETIONRAMWRITEDATAU2 (MICOMPLETIONRAMWRITEDATAU[2], MICOMPLETIONRAMWRITEDATAU_OUT[2]);
  buf B_MICOMPLETIONRAMWRITEDATAU20 (MICOMPLETIONRAMWRITEDATAU[20], MICOMPLETIONRAMWRITEDATAU_OUT[20]);
  buf B_MICOMPLETIONRAMWRITEDATAU21 (MICOMPLETIONRAMWRITEDATAU[21], MICOMPLETIONRAMWRITEDATAU_OUT[21]);
  buf B_MICOMPLETIONRAMWRITEDATAU22 (MICOMPLETIONRAMWRITEDATAU[22], MICOMPLETIONRAMWRITEDATAU_OUT[22]);
  buf B_MICOMPLETIONRAMWRITEDATAU23 (MICOMPLETIONRAMWRITEDATAU[23], MICOMPLETIONRAMWRITEDATAU_OUT[23]);
  buf B_MICOMPLETIONRAMWRITEDATAU24 (MICOMPLETIONRAMWRITEDATAU[24], MICOMPLETIONRAMWRITEDATAU_OUT[24]);
  buf B_MICOMPLETIONRAMWRITEDATAU25 (MICOMPLETIONRAMWRITEDATAU[25], MICOMPLETIONRAMWRITEDATAU_OUT[25]);
  buf B_MICOMPLETIONRAMWRITEDATAU26 (MICOMPLETIONRAMWRITEDATAU[26], MICOMPLETIONRAMWRITEDATAU_OUT[26]);
  buf B_MICOMPLETIONRAMWRITEDATAU27 (MICOMPLETIONRAMWRITEDATAU[27], MICOMPLETIONRAMWRITEDATAU_OUT[27]);
  buf B_MICOMPLETIONRAMWRITEDATAU28 (MICOMPLETIONRAMWRITEDATAU[28], MICOMPLETIONRAMWRITEDATAU_OUT[28]);
  buf B_MICOMPLETIONRAMWRITEDATAU29 (MICOMPLETIONRAMWRITEDATAU[29], MICOMPLETIONRAMWRITEDATAU_OUT[29]);
  buf B_MICOMPLETIONRAMWRITEDATAU3 (MICOMPLETIONRAMWRITEDATAU[3], MICOMPLETIONRAMWRITEDATAU_OUT[3]);
  buf B_MICOMPLETIONRAMWRITEDATAU30 (MICOMPLETIONRAMWRITEDATAU[30], MICOMPLETIONRAMWRITEDATAU_OUT[30]);
  buf B_MICOMPLETIONRAMWRITEDATAU31 (MICOMPLETIONRAMWRITEDATAU[31], MICOMPLETIONRAMWRITEDATAU_OUT[31]);
  buf B_MICOMPLETIONRAMWRITEDATAU32 (MICOMPLETIONRAMWRITEDATAU[32], MICOMPLETIONRAMWRITEDATAU_OUT[32]);
  buf B_MICOMPLETIONRAMWRITEDATAU33 (MICOMPLETIONRAMWRITEDATAU[33], MICOMPLETIONRAMWRITEDATAU_OUT[33]);
  buf B_MICOMPLETIONRAMWRITEDATAU34 (MICOMPLETIONRAMWRITEDATAU[34], MICOMPLETIONRAMWRITEDATAU_OUT[34]);
  buf B_MICOMPLETIONRAMWRITEDATAU35 (MICOMPLETIONRAMWRITEDATAU[35], MICOMPLETIONRAMWRITEDATAU_OUT[35]);
  buf B_MICOMPLETIONRAMWRITEDATAU36 (MICOMPLETIONRAMWRITEDATAU[36], MICOMPLETIONRAMWRITEDATAU_OUT[36]);
  buf B_MICOMPLETIONRAMWRITEDATAU37 (MICOMPLETIONRAMWRITEDATAU[37], MICOMPLETIONRAMWRITEDATAU_OUT[37]);
  buf B_MICOMPLETIONRAMWRITEDATAU38 (MICOMPLETIONRAMWRITEDATAU[38], MICOMPLETIONRAMWRITEDATAU_OUT[38]);
  buf B_MICOMPLETIONRAMWRITEDATAU39 (MICOMPLETIONRAMWRITEDATAU[39], MICOMPLETIONRAMWRITEDATAU_OUT[39]);
  buf B_MICOMPLETIONRAMWRITEDATAU4 (MICOMPLETIONRAMWRITEDATAU[4], MICOMPLETIONRAMWRITEDATAU_OUT[4]);
  buf B_MICOMPLETIONRAMWRITEDATAU40 (MICOMPLETIONRAMWRITEDATAU[40], MICOMPLETIONRAMWRITEDATAU_OUT[40]);
  buf B_MICOMPLETIONRAMWRITEDATAU41 (MICOMPLETIONRAMWRITEDATAU[41], MICOMPLETIONRAMWRITEDATAU_OUT[41]);
  buf B_MICOMPLETIONRAMWRITEDATAU42 (MICOMPLETIONRAMWRITEDATAU[42], MICOMPLETIONRAMWRITEDATAU_OUT[42]);
  buf B_MICOMPLETIONRAMWRITEDATAU43 (MICOMPLETIONRAMWRITEDATAU[43], MICOMPLETIONRAMWRITEDATAU_OUT[43]);
  buf B_MICOMPLETIONRAMWRITEDATAU44 (MICOMPLETIONRAMWRITEDATAU[44], MICOMPLETIONRAMWRITEDATAU_OUT[44]);
  buf B_MICOMPLETIONRAMWRITEDATAU45 (MICOMPLETIONRAMWRITEDATAU[45], MICOMPLETIONRAMWRITEDATAU_OUT[45]);
  buf B_MICOMPLETIONRAMWRITEDATAU46 (MICOMPLETIONRAMWRITEDATAU[46], MICOMPLETIONRAMWRITEDATAU_OUT[46]);
  buf B_MICOMPLETIONRAMWRITEDATAU47 (MICOMPLETIONRAMWRITEDATAU[47], MICOMPLETIONRAMWRITEDATAU_OUT[47]);
  buf B_MICOMPLETIONRAMWRITEDATAU48 (MICOMPLETIONRAMWRITEDATAU[48], MICOMPLETIONRAMWRITEDATAU_OUT[48]);
  buf B_MICOMPLETIONRAMWRITEDATAU49 (MICOMPLETIONRAMWRITEDATAU[49], MICOMPLETIONRAMWRITEDATAU_OUT[49]);
  buf B_MICOMPLETIONRAMWRITEDATAU5 (MICOMPLETIONRAMWRITEDATAU[5], MICOMPLETIONRAMWRITEDATAU_OUT[5]);
  buf B_MICOMPLETIONRAMWRITEDATAU50 (MICOMPLETIONRAMWRITEDATAU[50], MICOMPLETIONRAMWRITEDATAU_OUT[50]);
  buf B_MICOMPLETIONRAMWRITEDATAU51 (MICOMPLETIONRAMWRITEDATAU[51], MICOMPLETIONRAMWRITEDATAU_OUT[51]);
  buf B_MICOMPLETIONRAMWRITEDATAU52 (MICOMPLETIONRAMWRITEDATAU[52], MICOMPLETIONRAMWRITEDATAU_OUT[52]);
  buf B_MICOMPLETIONRAMWRITEDATAU53 (MICOMPLETIONRAMWRITEDATAU[53], MICOMPLETIONRAMWRITEDATAU_OUT[53]);
  buf B_MICOMPLETIONRAMWRITEDATAU54 (MICOMPLETIONRAMWRITEDATAU[54], MICOMPLETIONRAMWRITEDATAU_OUT[54]);
  buf B_MICOMPLETIONRAMWRITEDATAU55 (MICOMPLETIONRAMWRITEDATAU[55], MICOMPLETIONRAMWRITEDATAU_OUT[55]);
  buf B_MICOMPLETIONRAMWRITEDATAU56 (MICOMPLETIONRAMWRITEDATAU[56], MICOMPLETIONRAMWRITEDATAU_OUT[56]);
  buf B_MICOMPLETIONRAMWRITEDATAU57 (MICOMPLETIONRAMWRITEDATAU[57], MICOMPLETIONRAMWRITEDATAU_OUT[57]);
  buf B_MICOMPLETIONRAMWRITEDATAU58 (MICOMPLETIONRAMWRITEDATAU[58], MICOMPLETIONRAMWRITEDATAU_OUT[58]);
  buf B_MICOMPLETIONRAMWRITEDATAU59 (MICOMPLETIONRAMWRITEDATAU[59], MICOMPLETIONRAMWRITEDATAU_OUT[59]);
  buf B_MICOMPLETIONRAMWRITEDATAU6 (MICOMPLETIONRAMWRITEDATAU[6], MICOMPLETIONRAMWRITEDATAU_OUT[6]);
  buf B_MICOMPLETIONRAMWRITEDATAU60 (MICOMPLETIONRAMWRITEDATAU[60], MICOMPLETIONRAMWRITEDATAU_OUT[60]);
  buf B_MICOMPLETIONRAMWRITEDATAU61 (MICOMPLETIONRAMWRITEDATAU[61], MICOMPLETIONRAMWRITEDATAU_OUT[61]);
  buf B_MICOMPLETIONRAMWRITEDATAU62 (MICOMPLETIONRAMWRITEDATAU[62], MICOMPLETIONRAMWRITEDATAU_OUT[62]);
  buf B_MICOMPLETIONRAMWRITEDATAU63 (MICOMPLETIONRAMWRITEDATAU[63], MICOMPLETIONRAMWRITEDATAU_OUT[63]);
  buf B_MICOMPLETIONRAMWRITEDATAU64 (MICOMPLETIONRAMWRITEDATAU[64], MICOMPLETIONRAMWRITEDATAU_OUT[64]);
  buf B_MICOMPLETIONRAMWRITEDATAU65 (MICOMPLETIONRAMWRITEDATAU[65], MICOMPLETIONRAMWRITEDATAU_OUT[65]);
  buf B_MICOMPLETIONRAMWRITEDATAU66 (MICOMPLETIONRAMWRITEDATAU[66], MICOMPLETIONRAMWRITEDATAU_OUT[66]);
  buf B_MICOMPLETIONRAMWRITEDATAU67 (MICOMPLETIONRAMWRITEDATAU[67], MICOMPLETIONRAMWRITEDATAU_OUT[67]);
  buf B_MICOMPLETIONRAMWRITEDATAU68 (MICOMPLETIONRAMWRITEDATAU[68], MICOMPLETIONRAMWRITEDATAU_OUT[68]);
  buf B_MICOMPLETIONRAMWRITEDATAU69 (MICOMPLETIONRAMWRITEDATAU[69], MICOMPLETIONRAMWRITEDATAU_OUT[69]);
  buf B_MICOMPLETIONRAMWRITEDATAU7 (MICOMPLETIONRAMWRITEDATAU[7], MICOMPLETIONRAMWRITEDATAU_OUT[7]);
  buf B_MICOMPLETIONRAMWRITEDATAU70 (MICOMPLETIONRAMWRITEDATAU[70], MICOMPLETIONRAMWRITEDATAU_OUT[70]);
  buf B_MICOMPLETIONRAMWRITEDATAU71 (MICOMPLETIONRAMWRITEDATAU[71], MICOMPLETIONRAMWRITEDATAU_OUT[71]);
  buf B_MICOMPLETIONRAMWRITEDATAU8 (MICOMPLETIONRAMWRITEDATAU[8], MICOMPLETIONRAMWRITEDATAU_OUT[8]);
  buf B_MICOMPLETIONRAMWRITEDATAU9 (MICOMPLETIONRAMWRITEDATAU[9], MICOMPLETIONRAMWRITEDATAU_OUT[9]);
  buf B_MICOMPLETIONRAMWRITEENABLEL0 (MICOMPLETIONRAMWRITEENABLEL[0], MICOMPLETIONRAMWRITEENABLEL_OUT[0]);
  buf B_MICOMPLETIONRAMWRITEENABLEL1 (MICOMPLETIONRAMWRITEENABLEL[1], MICOMPLETIONRAMWRITEENABLEL_OUT[1]);
  buf B_MICOMPLETIONRAMWRITEENABLEL2 (MICOMPLETIONRAMWRITEENABLEL[2], MICOMPLETIONRAMWRITEENABLEL_OUT[2]);
  buf B_MICOMPLETIONRAMWRITEENABLEL3 (MICOMPLETIONRAMWRITEENABLEL[3], MICOMPLETIONRAMWRITEENABLEL_OUT[3]);
  buf B_MICOMPLETIONRAMWRITEENABLEU0 (MICOMPLETIONRAMWRITEENABLEU[0], MICOMPLETIONRAMWRITEENABLEU_OUT[0]);
  buf B_MICOMPLETIONRAMWRITEENABLEU1 (MICOMPLETIONRAMWRITEENABLEU[1], MICOMPLETIONRAMWRITEENABLEU_OUT[1]);
  buf B_MICOMPLETIONRAMWRITEENABLEU2 (MICOMPLETIONRAMWRITEENABLEU[2], MICOMPLETIONRAMWRITEENABLEU_OUT[2]);
  buf B_MICOMPLETIONRAMWRITEENABLEU3 (MICOMPLETIONRAMWRITEENABLEU[3], MICOMPLETIONRAMWRITEENABLEU_OUT[3]);
  buf B_MIREPLAYRAMADDRESS0 (MIREPLAYRAMADDRESS[0], MIREPLAYRAMADDRESS_OUT[0]);
  buf B_MIREPLAYRAMADDRESS1 (MIREPLAYRAMADDRESS[1], MIREPLAYRAMADDRESS_OUT[1]);
  buf B_MIREPLAYRAMADDRESS2 (MIREPLAYRAMADDRESS[2], MIREPLAYRAMADDRESS_OUT[2]);
  buf B_MIREPLAYRAMADDRESS3 (MIREPLAYRAMADDRESS[3], MIREPLAYRAMADDRESS_OUT[3]);
  buf B_MIREPLAYRAMADDRESS4 (MIREPLAYRAMADDRESS[4], MIREPLAYRAMADDRESS_OUT[4]);
  buf B_MIREPLAYRAMADDRESS5 (MIREPLAYRAMADDRESS[5], MIREPLAYRAMADDRESS_OUT[5]);
  buf B_MIREPLAYRAMADDRESS6 (MIREPLAYRAMADDRESS[6], MIREPLAYRAMADDRESS_OUT[6]);
  buf B_MIREPLAYRAMADDRESS7 (MIREPLAYRAMADDRESS[7], MIREPLAYRAMADDRESS_OUT[7]);
  buf B_MIREPLAYRAMADDRESS8 (MIREPLAYRAMADDRESS[8], MIREPLAYRAMADDRESS_OUT[8]);
  buf B_MIREPLAYRAMREADENABLE0 (MIREPLAYRAMREADENABLE[0], MIREPLAYRAMREADENABLE_OUT[0]);
  buf B_MIREPLAYRAMREADENABLE1 (MIREPLAYRAMREADENABLE[1], MIREPLAYRAMREADENABLE_OUT[1]);
  buf B_MIREPLAYRAMWRITEDATA0 (MIREPLAYRAMWRITEDATA[0], MIREPLAYRAMWRITEDATA_OUT[0]);
  buf B_MIREPLAYRAMWRITEDATA1 (MIREPLAYRAMWRITEDATA[1], MIREPLAYRAMWRITEDATA_OUT[1]);
  buf B_MIREPLAYRAMWRITEDATA10 (MIREPLAYRAMWRITEDATA[10], MIREPLAYRAMWRITEDATA_OUT[10]);
  buf B_MIREPLAYRAMWRITEDATA100 (MIREPLAYRAMWRITEDATA[100], MIREPLAYRAMWRITEDATA_OUT[100]);
  buf B_MIREPLAYRAMWRITEDATA101 (MIREPLAYRAMWRITEDATA[101], MIREPLAYRAMWRITEDATA_OUT[101]);
  buf B_MIREPLAYRAMWRITEDATA102 (MIREPLAYRAMWRITEDATA[102], MIREPLAYRAMWRITEDATA_OUT[102]);
  buf B_MIREPLAYRAMWRITEDATA103 (MIREPLAYRAMWRITEDATA[103], MIREPLAYRAMWRITEDATA_OUT[103]);
  buf B_MIREPLAYRAMWRITEDATA104 (MIREPLAYRAMWRITEDATA[104], MIREPLAYRAMWRITEDATA_OUT[104]);
  buf B_MIREPLAYRAMWRITEDATA105 (MIREPLAYRAMWRITEDATA[105], MIREPLAYRAMWRITEDATA_OUT[105]);
  buf B_MIREPLAYRAMWRITEDATA106 (MIREPLAYRAMWRITEDATA[106], MIREPLAYRAMWRITEDATA_OUT[106]);
  buf B_MIREPLAYRAMWRITEDATA107 (MIREPLAYRAMWRITEDATA[107], MIREPLAYRAMWRITEDATA_OUT[107]);
  buf B_MIREPLAYRAMWRITEDATA108 (MIREPLAYRAMWRITEDATA[108], MIREPLAYRAMWRITEDATA_OUT[108]);
  buf B_MIREPLAYRAMWRITEDATA109 (MIREPLAYRAMWRITEDATA[109], MIREPLAYRAMWRITEDATA_OUT[109]);
  buf B_MIREPLAYRAMWRITEDATA11 (MIREPLAYRAMWRITEDATA[11], MIREPLAYRAMWRITEDATA_OUT[11]);
  buf B_MIREPLAYRAMWRITEDATA110 (MIREPLAYRAMWRITEDATA[110], MIREPLAYRAMWRITEDATA_OUT[110]);
  buf B_MIREPLAYRAMWRITEDATA111 (MIREPLAYRAMWRITEDATA[111], MIREPLAYRAMWRITEDATA_OUT[111]);
  buf B_MIREPLAYRAMWRITEDATA112 (MIREPLAYRAMWRITEDATA[112], MIREPLAYRAMWRITEDATA_OUT[112]);
  buf B_MIREPLAYRAMWRITEDATA113 (MIREPLAYRAMWRITEDATA[113], MIREPLAYRAMWRITEDATA_OUT[113]);
  buf B_MIREPLAYRAMWRITEDATA114 (MIREPLAYRAMWRITEDATA[114], MIREPLAYRAMWRITEDATA_OUT[114]);
  buf B_MIREPLAYRAMWRITEDATA115 (MIREPLAYRAMWRITEDATA[115], MIREPLAYRAMWRITEDATA_OUT[115]);
  buf B_MIREPLAYRAMWRITEDATA116 (MIREPLAYRAMWRITEDATA[116], MIREPLAYRAMWRITEDATA_OUT[116]);
  buf B_MIREPLAYRAMWRITEDATA117 (MIREPLAYRAMWRITEDATA[117], MIREPLAYRAMWRITEDATA_OUT[117]);
  buf B_MIREPLAYRAMWRITEDATA118 (MIREPLAYRAMWRITEDATA[118], MIREPLAYRAMWRITEDATA_OUT[118]);
  buf B_MIREPLAYRAMWRITEDATA119 (MIREPLAYRAMWRITEDATA[119], MIREPLAYRAMWRITEDATA_OUT[119]);
  buf B_MIREPLAYRAMWRITEDATA12 (MIREPLAYRAMWRITEDATA[12], MIREPLAYRAMWRITEDATA_OUT[12]);
  buf B_MIREPLAYRAMWRITEDATA120 (MIREPLAYRAMWRITEDATA[120], MIREPLAYRAMWRITEDATA_OUT[120]);
  buf B_MIREPLAYRAMWRITEDATA121 (MIREPLAYRAMWRITEDATA[121], MIREPLAYRAMWRITEDATA_OUT[121]);
  buf B_MIREPLAYRAMWRITEDATA122 (MIREPLAYRAMWRITEDATA[122], MIREPLAYRAMWRITEDATA_OUT[122]);
  buf B_MIREPLAYRAMWRITEDATA123 (MIREPLAYRAMWRITEDATA[123], MIREPLAYRAMWRITEDATA_OUT[123]);
  buf B_MIREPLAYRAMWRITEDATA124 (MIREPLAYRAMWRITEDATA[124], MIREPLAYRAMWRITEDATA_OUT[124]);
  buf B_MIREPLAYRAMWRITEDATA125 (MIREPLAYRAMWRITEDATA[125], MIREPLAYRAMWRITEDATA_OUT[125]);
  buf B_MIREPLAYRAMWRITEDATA126 (MIREPLAYRAMWRITEDATA[126], MIREPLAYRAMWRITEDATA_OUT[126]);
  buf B_MIREPLAYRAMWRITEDATA127 (MIREPLAYRAMWRITEDATA[127], MIREPLAYRAMWRITEDATA_OUT[127]);
  buf B_MIREPLAYRAMWRITEDATA128 (MIREPLAYRAMWRITEDATA[128], MIREPLAYRAMWRITEDATA_OUT[128]);
  buf B_MIREPLAYRAMWRITEDATA129 (MIREPLAYRAMWRITEDATA[129], MIREPLAYRAMWRITEDATA_OUT[129]);
  buf B_MIREPLAYRAMWRITEDATA13 (MIREPLAYRAMWRITEDATA[13], MIREPLAYRAMWRITEDATA_OUT[13]);
  buf B_MIREPLAYRAMWRITEDATA130 (MIREPLAYRAMWRITEDATA[130], MIREPLAYRAMWRITEDATA_OUT[130]);
  buf B_MIREPLAYRAMWRITEDATA131 (MIREPLAYRAMWRITEDATA[131], MIREPLAYRAMWRITEDATA_OUT[131]);
  buf B_MIREPLAYRAMWRITEDATA132 (MIREPLAYRAMWRITEDATA[132], MIREPLAYRAMWRITEDATA_OUT[132]);
  buf B_MIREPLAYRAMWRITEDATA133 (MIREPLAYRAMWRITEDATA[133], MIREPLAYRAMWRITEDATA_OUT[133]);
  buf B_MIREPLAYRAMWRITEDATA134 (MIREPLAYRAMWRITEDATA[134], MIREPLAYRAMWRITEDATA_OUT[134]);
  buf B_MIREPLAYRAMWRITEDATA135 (MIREPLAYRAMWRITEDATA[135], MIREPLAYRAMWRITEDATA_OUT[135]);
  buf B_MIREPLAYRAMWRITEDATA136 (MIREPLAYRAMWRITEDATA[136], MIREPLAYRAMWRITEDATA_OUT[136]);
  buf B_MIREPLAYRAMWRITEDATA137 (MIREPLAYRAMWRITEDATA[137], MIREPLAYRAMWRITEDATA_OUT[137]);
  buf B_MIREPLAYRAMWRITEDATA138 (MIREPLAYRAMWRITEDATA[138], MIREPLAYRAMWRITEDATA_OUT[138]);
  buf B_MIREPLAYRAMWRITEDATA139 (MIREPLAYRAMWRITEDATA[139], MIREPLAYRAMWRITEDATA_OUT[139]);
  buf B_MIREPLAYRAMWRITEDATA14 (MIREPLAYRAMWRITEDATA[14], MIREPLAYRAMWRITEDATA_OUT[14]);
  buf B_MIREPLAYRAMWRITEDATA140 (MIREPLAYRAMWRITEDATA[140], MIREPLAYRAMWRITEDATA_OUT[140]);
  buf B_MIREPLAYRAMWRITEDATA141 (MIREPLAYRAMWRITEDATA[141], MIREPLAYRAMWRITEDATA_OUT[141]);
  buf B_MIREPLAYRAMWRITEDATA142 (MIREPLAYRAMWRITEDATA[142], MIREPLAYRAMWRITEDATA_OUT[142]);
  buf B_MIREPLAYRAMWRITEDATA143 (MIREPLAYRAMWRITEDATA[143], MIREPLAYRAMWRITEDATA_OUT[143]);
  buf B_MIREPLAYRAMWRITEDATA15 (MIREPLAYRAMWRITEDATA[15], MIREPLAYRAMWRITEDATA_OUT[15]);
  buf B_MIREPLAYRAMWRITEDATA16 (MIREPLAYRAMWRITEDATA[16], MIREPLAYRAMWRITEDATA_OUT[16]);
  buf B_MIREPLAYRAMWRITEDATA17 (MIREPLAYRAMWRITEDATA[17], MIREPLAYRAMWRITEDATA_OUT[17]);
  buf B_MIREPLAYRAMWRITEDATA18 (MIREPLAYRAMWRITEDATA[18], MIREPLAYRAMWRITEDATA_OUT[18]);
  buf B_MIREPLAYRAMWRITEDATA19 (MIREPLAYRAMWRITEDATA[19], MIREPLAYRAMWRITEDATA_OUT[19]);
  buf B_MIREPLAYRAMWRITEDATA2 (MIREPLAYRAMWRITEDATA[2], MIREPLAYRAMWRITEDATA_OUT[2]);
  buf B_MIREPLAYRAMWRITEDATA20 (MIREPLAYRAMWRITEDATA[20], MIREPLAYRAMWRITEDATA_OUT[20]);
  buf B_MIREPLAYRAMWRITEDATA21 (MIREPLAYRAMWRITEDATA[21], MIREPLAYRAMWRITEDATA_OUT[21]);
  buf B_MIREPLAYRAMWRITEDATA22 (MIREPLAYRAMWRITEDATA[22], MIREPLAYRAMWRITEDATA_OUT[22]);
  buf B_MIREPLAYRAMWRITEDATA23 (MIREPLAYRAMWRITEDATA[23], MIREPLAYRAMWRITEDATA_OUT[23]);
  buf B_MIREPLAYRAMWRITEDATA24 (MIREPLAYRAMWRITEDATA[24], MIREPLAYRAMWRITEDATA_OUT[24]);
  buf B_MIREPLAYRAMWRITEDATA25 (MIREPLAYRAMWRITEDATA[25], MIREPLAYRAMWRITEDATA_OUT[25]);
  buf B_MIREPLAYRAMWRITEDATA26 (MIREPLAYRAMWRITEDATA[26], MIREPLAYRAMWRITEDATA_OUT[26]);
  buf B_MIREPLAYRAMWRITEDATA27 (MIREPLAYRAMWRITEDATA[27], MIREPLAYRAMWRITEDATA_OUT[27]);
  buf B_MIREPLAYRAMWRITEDATA28 (MIREPLAYRAMWRITEDATA[28], MIREPLAYRAMWRITEDATA_OUT[28]);
  buf B_MIREPLAYRAMWRITEDATA29 (MIREPLAYRAMWRITEDATA[29], MIREPLAYRAMWRITEDATA_OUT[29]);
  buf B_MIREPLAYRAMWRITEDATA3 (MIREPLAYRAMWRITEDATA[3], MIREPLAYRAMWRITEDATA_OUT[3]);
  buf B_MIREPLAYRAMWRITEDATA30 (MIREPLAYRAMWRITEDATA[30], MIREPLAYRAMWRITEDATA_OUT[30]);
  buf B_MIREPLAYRAMWRITEDATA31 (MIREPLAYRAMWRITEDATA[31], MIREPLAYRAMWRITEDATA_OUT[31]);
  buf B_MIREPLAYRAMWRITEDATA32 (MIREPLAYRAMWRITEDATA[32], MIREPLAYRAMWRITEDATA_OUT[32]);
  buf B_MIREPLAYRAMWRITEDATA33 (MIREPLAYRAMWRITEDATA[33], MIREPLAYRAMWRITEDATA_OUT[33]);
  buf B_MIREPLAYRAMWRITEDATA34 (MIREPLAYRAMWRITEDATA[34], MIREPLAYRAMWRITEDATA_OUT[34]);
  buf B_MIREPLAYRAMWRITEDATA35 (MIREPLAYRAMWRITEDATA[35], MIREPLAYRAMWRITEDATA_OUT[35]);
  buf B_MIREPLAYRAMWRITEDATA36 (MIREPLAYRAMWRITEDATA[36], MIREPLAYRAMWRITEDATA_OUT[36]);
  buf B_MIREPLAYRAMWRITEDATA37 (MIREPLAYRAMWRITEDATA[37], MIREPLAYRAMWRITEDATA_OUT[37]);
  buf B_MIREPLAYRAMWRITEDATA38 (MIREPLAYRAMWRITEDATA[38], MIREPLAYRAMWRITEDATA_OUT[38]);
  buf B_MIREPLAYRAMWRITEDATA39 (MIREPLAYRAMWRITEDATA[39], MIREPLAYRAMWRITEDATA_OUT[39]);
  buf B_MIREPLAYRAMWRITEDATA4 (MIREPLAYRAMWRITEDATA[4], MIREPLAYRAMWRITEDATA_OUT[4]);
  buf B_MIREPLAYRAMWRITEDATA40 (MIREPLAYRAMWRITEDATA[40], MIREPLAYRAMWRITEDATA_OUT[40]);
  buf B_MIREPLAYRAMWRITEDATA41 (MIREPLAYRAMWRITEDATA[41], MIREPLAYRAMWRITEDATA_OUT[41]);
  buf B_MIREPLAYRAMWRITEDATA42 (MIREPLAYRAMWRITEDATA[42], MIREPLAYRAMWRITEDATA_OUT[42]);
  buf B_MIREPLAYRAMWRITEDATA43 (MIREPLAYRAMWRITEDATA[43], MIREPLAYRAMWRITEDATA_OUT[43]);
  buf B_MIREPLAYRAMWRITEDATA44 (MIREPLAYRAMWRITEDATA[44], MIREPLAYRAMWRITEDATA_OUT[44]);
  buf B_MIREPLAYRAMWRITEDATA45 (MIREPLAYRAMWRITEDATA[45], MIREPLAYRAMWRITEDATA_OUT[45]);
  buf B_MIREPLAYRAMWRITEDATA46 (MIREPLAYRAMWRITEDATA[46], MIREPLAYRAMWRITEDATA_OUT[46]);
  buf B_MIREPLAYRAMWRITEDATA47 (MIREPLAYRAMWRITEDATA[47], MIREPLAYRAMWRITEDATA_OUT[47]);
  buf B_MIREPLAYRAMWRITEDATA48 (MIREPLAYRAMWRITEDATA[48], MIREPLAYRAMWRITEDATA_OUT[48]);
  buf B_MIREPLAYRAMWRITEDATA49 (MIREPLAYRAMWRITEDATA[49], MIREPLAYRAMWRITEDATA_OUT[49]);
  buf B_MIREPLAYRAMWRITEDATA5 (MIREPLAYRAMWRITEDATA[5], MIREPLAYRAMWRITEDATA_OUT[5]);
  buf B_MIREPLAYRAMWRITEDATA50 (MIREPLAYRAMWRITEDATA[50], MIREPLAYRAMWRITEDATA_OUT[50]);
  buf B_MIREPLAYRAMWRITEDATA51 (MIREPLAYRAMWRITEDATA[51], MIREPLAYRAMWRITEDATA_OUT[51]);
  buf B_MIREPLAYRAMWRITEDATA52 (MIREPLAYRAMWRITEDATA[52], MIREPLAYRAMWRITEDATA_OUT[52]);
  buf B_MIREPLAYRAMWRITEDATA53 (MIREPLAYRAMWRITEDATA[53], MIREPLAYRAMWRITEDATA_OUT[53]);
  buf B_MIREPLAYRAMWRITEDATA54 (MIREPLAYRAMWRITEDATA[54], MIREPLAYRAMWRITEDATA_OUT[54]);
  buf B_MIREPLAYRAMWRITEDATA55 (MIREPLAYRAMWRITEDATA[55], MIREPLAYRAMWRITEDATA_OUT[55]);
  buf B_MIREPLAYRAMWRITEDATA56 (MIREPLAYRAMWRITEDATA[56], MIREPLAYRAMWRITEDATA_OUT[56]);
  buf B_MIREPLAYRAMWRITEDATA57 (MIREPLAYRAMWRITEDATA[57], MIREPLAYRAMWRITEDATA_OUT[57]);
  buf B_MIREPLAYRAMWRITEDATA58 (MIREPLAYRAMWRITEDATA[58], MIREPLAYRAMWRITEDATA_OUT[58]);
  buf B_MIREPLAYRAMWRITEDATA59 (MIREPLAYRAMWRITEDATA[59], MIREPLAYRAMWRITEDATA_OUT[59]);
  buf B_MIREPLAYRAMWRITEDATA6 (MIREPLAYRAMWRITEDATA[6], MIREPLAYRAMWRITEDATA_OUT[6]);
  buf B_MIREPLAYRAMWRITEDATA60 (MIREPLAYRAMWRITEDATA[60], MIREPLAYRAMWRITEDATA_OUT[60]);
  buf B_MIREPLAYRAMWRITEDATA61 (MIREPLAYRAMWRITEDATA[61], MIREPLAYRAMWRITEDATA_OUT[61]);
  buf B_MIREPLAYRAMWRITEDATA62 (MIREPLAYRAMWRITEDATA[62], MIREPLAYRAMWRITEDATA_OUT[62]);
  buf B_MIREPLAYRAMWRITEDATA63 (MIREPLAYRAMWRITEDATA[63], MIREPLAYRAMWRITEDATA_OUT[63]);
  buf B_MIREPLAYRAMWRITEDATA64 (MIREPLAYRAMWRITEDATA[64], MIREPLAYRAMWRITEDATA_OUT[64]);
  buf B_MIREPLAYRAMWRITEDATA65 (MIREPLAYRAMWRITEDATA[65], MIREPLAYRAMWRITEDATA_OUT[65]);
  buf B_MIREPLAYRAMWRITEDATA66 (MIREPLAYRAMWRITEDATA[66], MIREPLAYRAMWRITEDATA_OUT[66]);
  buf B_MIREPLAYRAMWRITEDATA67 (MIREPLAYRAMWRITEDATA[67], MIREPLAYRAMWRITEDATA_OUT[67]);
  buf B_MIREPLAYRAMWRITEDATA68 (MIREPLAYRAMWRITEDATA[68], MIREPLAYRAMWRITEDATA_OUT[68]);
  buf B_MIREPLAYRAMWRITEDATA69 (MIREPLAYRAMWRITEDATA[69], MIREPLAYRAMWRITEDATA_OUT[69]);
  buf B_MIREPLAYRAMWRITEDATA7 (MIREPLAYRAMWRITEDATA[7], MIREPLAYRAMWRITEDATA_OUT[7]);
  buf B_MIREPLAYRAMWRITEDATA70 (MIREPLAYRAMWRITEDATA[70], MIREPLAYRAMWRITEDATA_OUT[70]);
  buf B_MIREPLAYRAMWRITEDATA71 (MIREPLAYRAMWRITEDATA[71], MIREPLAYRAMWRITEDATA_OUT[71]);
  buf B_MIREPLAYRAMWRITEDATA72 (MIREPLAYRAMWRITEDATA[72], MIREPLAYRAMWRITEDATA_OUT[72]);
  buf B_MIREPLAYRAMWRITEDATA73 (MIREPLAYRAMWRITEDATA[73], MIREPLAYRAMWRITEDATA_OUT[73]);
  buf B_MIREPLAYRAMWRITEDATA74 (MIREPLAYRAMWRITEDATA[74], MIREPLAYRAMWRITEDATA_OUT[74]);
  buf B_MIREPLAYRAMWRITEDATA75 (MIREPLAYRAMWRITEDATA[75], MIREPLAYRAMWRITEDATA_OUT[75]);
  buf B_MIREPLAYRAMWRITEDATA76 (MIREPLAYRAMWRITEDATA[76], MIREPLAYRAMWRITEDATA_OUT[76]);
  buf B_MIREPLAYRAMWRITEDATA77 (MIREPLAYRAMWRITEDATA[77], MIREPLAYRAMWRITEDATA_OUT[77]);
  buf B_MIREPLAYRAMWRITEDATA78 (MIREPLAYRAMWRITEDATA[78], MIREPLAYRAMWRITEDATA_OUT[78]);
  buf B_MIREPLAYRAMWRITEDATA79 (MIREPLAYRAMWRITEDATA[79], MIREPLAYRAMWRITEDATA_OUT[79]);
  buf B_MIREPLAYRAMWRITEDATA8 (MIREPLAYRAMWRITEDATA[8], MIREPLAYRAMWRITEDATA_OUT[8]);
  buf B_MIREPLAYRAMWRITEDATA80 (MIREPLAYRAMWRITEDATA[80], MIREPLAYRAMWRITEDATA_OUT[80]);
  buf B_MIREPLAYRAMWRITEDATA81 (MIREPLAYRAMWRITEDATA[81], MIREPLAYRAMWRITEDATA_OUT[81]);
  buf B_MIREPLAYRAMWRITEDATA82 (MIREPLAYRAMWRITEDATA[82], MIREPLAYRAMWRITEDATA_OUT[82]);
  buf B_MIREPLAYRAMWRITEDATA83 (MIREPLAYRAMWRITEDATA[83], MIREPLAYRAMWRITEDATA_OUT[83]);
  buf B_MIREPLAYRAMWRITEDATA84 (MIREPLAYRAMWRITEDATA[84], MIREPLAYRAMWRITEDATA_OUT[84]);
  buf B_MIREPLAYRAMWRITEDATA85 (MIREPLAYRAMWRITEDATA[85], MIREPLAYRAMWRITEDATA_OUT[85]);
  buf B_MIREPLAYRAMWRITEDATA86 (MIREPLAYRAMWRITEDATA[86], MIREPLAYRAMWRITEDATA_OUT[86]);
  buf B_MIREPLAYRAMWRITEDATA87 (MIREPLAYRAMWRITEDATA[87], MIREPLAYRAMWRITEDATA_OUT[87]);
  buf B_MIREPLAYRAMWRITEDATA88 (MIREPLAYRAMWRITEDATA[88], MIREPLAYRAMWRITEDATA_OUT[88]);
  buf B_MIREPLAYRAMWRITEDATA89 (MIREPLAYRAMWRITEDATA[89], MIREPLAYRAMWRITEDATA_OUT[89]);
  buf B_MIREPLAYRAMWRITEDATA9 (MIREPLAYRAMWRITEDATA[9], MIREPLAYRAMWRITEDATA_OUT[9]);
  buf B_MIREPLAYRAMWRITEDATA90 (MIREPLAYRAMWRITEDATA[90], MIREPLAYRAMWRITEDATA_OUT[90]);
  buf B_MIREPLAYRAMWRITEDATA91 (MIREPLAYRAMWRITEDATA[91], MIREPLAYRAMWRITEDATA_OUT[91]);
  buf B_MIREPLAYRAMWRITEDATA92 (MIREPLAYRAMWRITEDATA[92], MIREPLAYRAMWRITEDATA_OUT[92]);
  buf B_MIREPLAYRAMWRITEDATA93 (MIREPLAYRAMWRITEDATA[93], MIREPLAYRAMWRITEDATA_OUT[93]);
  buf B_MIREPLAYRAMWRITEDATA94 (MIREPLAYRAMWRITEDATA[94], MIREPLAYRAMWRITEDATA_OUT[94]);
  buf B_MIREPLAYRAMWRITEDATA95 (MIREPLAYRAMWRITEDATA[95], MIREPLAYRAMWRITEDATA_OUT[95]);
  buf B_MIREPLAYRAMWRITEDATA96 (MIREPLAYRAMWRITEDATA[96], MIREPLAYRAMWRITEDATA_OUT[96]);
  buf B_MIREPLAYRAMWRITEDATA97 (MIREPLAYRAMWRITEDATA[97], MIREPLAYRAMWRITEDATA_OUT[97]);
  buf B_MIREPLAYRAMWRITEDATA98 (MIREPLAYRAMWRITEDATA[98], MIREPLAYRAMWRITEDATA_OUT[98]);
  buf B_MIREPLAYRAMWRITEDATA99 (MIREPLAYRAMWRITEDATA[99], MIREPLAYRAMWRITEDATA_OUT[99]);
  buf B_MIREPLAYRAMWRITEENABLE0 (MIREPLAYRAMWRITEENABLE[0], MIREPLAYRAMWRITEENABLE_OUT[0]);
  buf B_MIREPLAYRAMWRITEENABLE1 (MIREPLAYRAMWRITEENABLE[1], MIREPLAYRAMWRITEENABLE_OUT[1]);
  buf B_MIREQUESTRAMREADADDRESSA0 (MIREQUESTRAMREADADDRESSA[0], MIREQUESTRAMREADADDRESSA_OUT[0]);
  buf B_MIREQUESTRAMREADADDRESSA1 (MIREQUESTRAMREADADDRESSA[1], MIREQUESTRAMREADADDRESSA_OUT[1]);
  buf B_MIREQUESTRAMREADADDRESSA2 (MIREQUESTRAMREADADDRESSA[2], MIREQUESTRAMREADADDRESSA_OUT[2]);
  buf B_MIREQUESTRAMREADADDRESSA3 (MIREQUESTRAMREADADDRESSA[3], MIREQUESTRAMREADADDRESSA_OUT[3]);
  buf B_MIREQUESTRAMREADADDRESSA4 (MIREQUESTRAMREADADDRESSA[4], MIREQUESTRAMREADADDRESSA_OUT[4]);
  buf B_MIREQUESTRAMREADADDRESSA5 (MIREQUESTRAMREADADDRESSA[5], MIREQUESTRAMREADADDRESSA_OUT[5]);
  buf B_MIREQUESTRAMREADADDRESSA6 (MIREQUESTRAMREADADDRESSA[6], MIREQUESTRAMREADADDRESSA_OUT[6]);
  buf B_MIREQUESTRAMREADADDRESSA7 (MIREQUESTRAMREADADDRESSA[7], MIREQUESTRAMREADADDRESSA_OUT[7]);
  buf B_MIREQUESTRAMREADADDRESSA8 (MIREQUESTRAMREADADDRESSA[8], MIREQUESTRAMREADADDRESSA_OUT[8]);
  buf B_MIREQUESTRAMREADADDRESSB0 (MIREQUESTRAMREADADDRESSB[0], MIREQUESTRAMREADADDRESSB_OUT[0]);
  buf B_MIREQUESTRAMREADADDRESSB1 (MIREQUESTRAMREADADDRESSB[1], MIREQUESTRAMREADADDRESSB_OUT[1]);
  buf B_MIREQUESTRAMREADADDRESSB2 (MIREQUESTRAMREADADDRESSB[2], MIREQUESTRAMREADADDRESSB_OUT[2]);
  buf B_MIREQUESTRAMREADADDRESSB3 (MIREQUESTRAMREADADDRESSB[3], MIREQUESTRAMREADADDRESSB_OUT[3]);
  buf B_MIREQUESTRAMREADADDRESSB4 (MIREQUESTRAMREADADDRESSB[4], MIREQUESTRAMREADADDRESSB_OUT[4]);
  buf B_MIREQUESTRAMREADADDRESSB5 (MIREQUESTRAMREADADDRESSB[5], MIREQUESTRAMREADADDRESSB_OUT[5]);
  buf B_MIREQUESTRAMREADADDRESSB6 (MIREQUESTRAMREADADDRESSB[6], MIREQUESTRAMREADADDRESSB_OUT[6]);
  buf B_MIREQUESTRAMREADADDRESSB7 (MIREQUESTRAMREADADDRESSB[7], MIREQUESTRAMREADADDRESSB_OUT[7]);
  buf B_MIREQUESTRAMREADADDRESSB8 (MIREQUESTRAMREADADDRESSB[8], MIREQUESTRAMREADADDRESSB_OUT[8]);
  buf B_MIREQUESTRAMREADENABLE0 (MIREQUESTRAMREADENABLE[0], MIREQUESTRAMREADENABLE_OUT[0]);
  buf B_MIREQUESTRAMREADENABLE1 (MIREQUESTRAMREADENABLE[1], MIREQUESTRAMREADENABLE_OUT[1]);
  buf B_MIREQUESTRAMREADENABLE2 (MIREQUESTRAMREADENABLE[2], MIREQUESTRAMREADENABLE_OUT[2]);
  buf B_MIREQUESTRAMREADENABLE3 (MIREQUESTRAMREADENABLE[3], MIREQUESTRAMREADENABLE_OUT[3]);
  buf B_MIREQUESTRAMWRITEADDRESSA0 (MIREQUESTRAMWRITEADDRESSA[0], MIREQUESTRAMWRITEADDRESSA_OUT[0]);
  buf B_MIREQUESTRAMWRITEADDRESSA1 (MIREQUESTRAMWRITEADDRESSA[1], MIREQUESTRAMWRITEADDRESSA_OUT[1]);
  buf B_MIREQUESTRAMWRITEADDRESSA2 (MIREQUESTRAMWRITEADDRESSA[2], MIREQUESTRAMWRITEADDRESSA_OUT[2]);
  buf B_MIREQUESTRAMWRITEADDRESSA3 (MIREQUESTRAMWRITEADDRESSA[3], MIREQUESTRAMWRITEADDRESSA_OUT[3]);
  buf B_MIREQUESTRAMWRITEADDRESSA4 (MIREQUESTRAMWRITEADDRESSA[4], MIREQUESTRAMWRITEADDRESSA_OUT[4]);
  buf B_MIREQUESTRAMWRITEADDRESSA5 (MIREQUESTRAMWRITEADDRESSA[5], MIREQUESTRAMWRITEADDRESSA_OUT[5]);
  buf B_MIREQUESTRAMWRITEADDRESSA6 (MIREQUESTRAMWRITEADDRESSA[6], MIREQUESTRAMWRITEADDRESSA_OUT[6]);
  buf B_MIREQUESTRAMWRITEADDRESSA7 (MIREQUESTRAMWRITEADDRESSA[7], MIREQUESTRAMWRITEADDRESSA_OUT[7]);
  buf B_MIREQUESTRAMWRITEADDRESSA8 (MIREQUESTRAMWRITEADDRESSA[8], MIREQUESTRAMWRITEADDRESSA_OUT[8]);
  buf B_MIREQUESTRAMWRITEADDRESSB0 (MIREQUESTRAMWRITEADDRESSB[0], MIREQUESTRAMWRITEADDRESSB_OUT[0]);
  buf B_MIREQUESTRAMWRITEADDRESSB1 (MIREQUESTRAMWRITEADDRESSB[1], MIREQUESTRAMWRITEADDRESSB_OUT[1]);
  buf B_MIREQUESTRAMWRITEADDRESSB2 (MIREQUESTRAMWRITEADDRESSB[2], MIREQUESTRAMWRITEADDRESSB_OUT[2]);
  buf B_MIREQUESTRAMWRITEADDRESSB3 (MIREQUESTRAMWRITEADDRESSB[3], MIREQUESTRAMWRITEADDRESSB_OUT[3]);
  buf B_MIREQUESTRAMWRITEADDRESSB4 (MIREQUESTRAMWRITEADDRESSB[4], MIREQUESTRAMWRITEADDRESSB_OUT[4]);
  buf B_MIREQUESTRAMWRITEADDRESSB5 (MIREQUESTRAMWRITEADDRESSB[5], MIREQUESTRAMWRITEADDRESSB_OUT[5]);
  buf B_MIREQUESTRAMWRITEADDRESSB6 (MIREQUESTRAMWRITEADDRESSB[6], MIREQUESTRAMWRITEADDRESSB_OUT[6]);
  buf B_MIREQUESTRAMWRITEADDRESSB7 (MIREQUESTRAMWRITEADDRESSB[7], MIREQUESTRAMWRITEADDRESSB_OUT[7]);
  buf B_MIREQUESTRAMWRITEADDRESSB8 (MIREQUESTRAMWRITEADDRESSB[8], MIREQUESTRAMWRITEADDRESSB_OUT[8]);
  buf B_MIREQUESTRAMWRITEDATA0 (MIREQUESTRAMWRITEDATA[0], MIREQUESTRAMWRITEDATA_OUT[0]);
  buf B_MIREQUESTRAMWRITEDATA1 (MIREQUESTRAMWRITEDATA[1], MIREQUESTRAMWRITEDATA_OUT[1]);
  buf B_MIREQUESTRAMWRITEDATA10 (MIREQUESTRAMWRITEDATA[10], MIREQUESTRAMWRITEDATA_OUT[10]);
  buf B_MIREQUESTRAMWRITEDATA100 (MIREQUESTRAMWRITEDATA[100], MIREQUESTRAMWRITEDATA_OUT[100]);
  buf B_MIREQUESTRAMWRITEDATA101 (MIREQUESTRAMWRITEDATA[101], MIREQUESTRAMWRITEDATA_OUT[101]);
  buf B_MIREQUESTRAMWRITEDATA102 (MIREQUESTRAMWRITEDATA[102], MIREQUESTRAMWRITEDATA_OUT[102]);
  buf B_MIREQUESTRAMWRITEDATA103 (MIREQUESTRAMWRITEDATA[103], MIREQUESTRAMWRITEDATA_OUT[103]);
  buf B_MIREQUESTRAMWRITEDATA104 (MIREQUESTRAMWRITEDATA[104], MIREQUESTRAMWRITEDATA_OUT[104]);
  buf B_MIREQUESTRAMWRITEDATA105 (MIREQUESTRAMWRITEDATA[105], MIREQUESTRAMWRITEDATA_OUT[105]);
  buf B_MIREQUESTRAMWRITEDATA106 (MIREQUESTRAMWRITEDATA[106], MIREQUESTRAMWRITEDATA_OUT[106]);
  buf B_MIREQUESTRAMWRITEDATA107 (MIREQUESTRAMWRITEDATA[107], MIREQUESTRAMWRITEDATA_OUT[107]);
  buf B_MIREQUESTRAMWRITEDATA108 (MIREQUESTRAMWRITEDATA[108], MIREQUESTRAMWRITEDATA_OUT[108]);
  buf B_MIREQUESTRAMWRITEDATA109 (MIREQUESTRAMWRITEDATA[109], MIREQUESTRAMWRITEDATA_OUT[109]);
  buf B_MIREQUESTRAMWRITEDATA11 (MIREQUESTRAMWRITEDATA[11], MIREQUESTRAMWRITEDATA_OUT[11]);
  buf B_MIREQUESTRAMWRITEDATA110 (MIREQUESTRAMWRITEDATA[110], MIREQUESTRAMWRITEDATA_OUT[110]);
  buf B_MIREQUESTRAMWRITEDATA111 (MIREQUESTRAMWRITEDATA[111], MIREQUESTRAMWRITEDATA_OUT[111]);
  buf B_MIREQUESTRAMWRITEDATA112 (MIREQUESTRAMWRITEDATA[112], MIREQUESTRAMWRITEDATA_OUT[112]);
  buf B_MIREQUESTRAMWRITEDATA113 (MIREQUESTRAMWRITEDATA[113], MIREQUESTRAMWRITEDATA_OUT[113]);
  buf B_MIREQUESTRAMWRITEDATA114 (MIREQUESTRAMWRITEDATA[114], MIREQUESTRAMWRITEDATA_OUT[114]);
  buf B_MIREQUESTRAMWRITEDATA115 (MIREQUESTRAMWRITEDATA[115], MIREQUESTRAMWRITEDATA_OUT[115]);
  buf B_MIREQUESTRAMWRITEDATA116 (MIREQUESTRAMWRITEDATA[116], MIREQUESTRAMWRITEDATA_OUT[116]);
  buf B_MIREQUESTRAMWRITEDATA117 (MIREQUESTRAMWRITEDATA[117], MIREQUESTRAMWRITEDATA_OUT[117]);
  buf B_MIREQUESTRAMWRITEDATA118 (MIREQUESTRAMWRITEDATA[118], MIREQUESTRAMWRITEDATA_OUT[118]);
  buf B_MIREQUESTRAMWRITEDATA119 (MIREQUESTRAMWRITEDATA[119], MIREQUESTRAMWRITEDATA_OUT[119]);
  buf B_MIREQUESTRAMWRITEDATA12 (MIREQUESTRAMWRITEDATA[12], MIREQUESTRAMWRITEDATA_OUT[12]);
  buf B_MIREQUESTRAMWRITEDATA120 (MIREQUESTRAMWRITEDATA[120], MIREQUESTRAMWRITEDATA_OUT[120]);
  buf B_MIREQUESTRAMWRITEDATA121 (MIREQUESTRAMWRITEDATA[121], MIREQUESTRAMWRITEDATA_OUT[121]);
  buf B_MIREQUESTRAMWRITEDATA122 (MIREQUESTRAMWRITEDATA[122], MIREQUESTRAMWRITEDATA_OUT[122]);
  buf B_MIREQUESTRAMWRITEDATA123 (MIREQUESTRAMWRITEDATA[123], MIREQUESTRAMWRITEDATA_OUT[123]);
  buf B_MIREQUESTRAMWRITEDATA124 (MIREQUESTRAMWRITEDATA[124], MIREQUESTRAMWRITEDATA_OUT[124]);
  buf B_MIREQUESTRAMWRITEDATA125 (MIREQUESTRAMWRITEDATA[125], MIREQUESTRAMWRITEDATA_OUT[125]);
  buf B_MIREQUESTRAMWRITEDATA126 (MIREQUESTRAMWRITEDATA[126], MIREQUESTRAMWRITEDATA_OUT[126]);
  buf B_MIREQUESTRAMWRITEDATA127 (MIREQUESTRAMWRITEDATA[127], MIREQUESTRAMWRITEDATA_OUT[127]);
  buf B_MIREQUESTRAMWRITEDATA128 (MIREQUESTRAMWRITEDATA[128], MIREQUESTRAMWRITEDATA_OUT[128]);
  buf B_MIREQUESTRAMWRITEDATA129 (MIREQUESTRAMWRITEDATA[129], MIREQUESTRAMWRITEDATA_OUT[129]);
  buf B_MIREQUESTRAMWRITEDATA13 (MIREQUESTRAMWRITEDATA[13], MIREQUESTRAMWRITEDATA_OUT[13]);
  buf B_MIREQUESTRAMWRITEDATA130 (MIREQUESTRAMWRITEDATA[130], MIREQUESTRAMWRITEDATA_OUT[130]);
  buf B_MIREQUESTRAMWRITEDATA131 (MIREQUESTRAMWRITEDATA[131], MIREQUESTRAMWRITEDATA_OUT[131]);
  buf B_MIREQUESTRAMWRITEDATA132 (MIREQUESTRAMWRITEDATA[132], MIREQUESTRAMWRITEDATA_OUT[132]);
  buf B_MIREQUESTRAMWRITEDATA133 (MIREQUESTRAMWRITEDATA[133], MIREQUESTRAMWRITEDATA_OUT[133]);
  buf B_MIREQUESTRAMWRITEDATA134 (MIREQUESTRAMWRITEDATA[134], MIREQUESTRAMWRITEDATA_OUT[134]);
  buf B_MIREQUESTRAMWRITEDATA135 (MIREQUESTRAMWRITEDATA[135], MIREQUESTRAMWRITEDATA_OUT[135]);
  buf B_MIREQUESTRAMWRITEDATA136 (MIREQUESTRAMWRITEDATA[136], MIREQUESTRAMWRITEDATA_OUT[136]);
  buf B_MIREQUESTRAMWRITEDATA137 (MIREQUESTRAMWRITEDATA[137], MIREQUESTRAMWRITEDATA_OUT[137]);
  buf B_MIREQUESTRAMWRITEDATA138 (MIREQUESTRAMWRITEDATA[138], MIREQUESTRAMWRITEDATA_OUT[138]);
  buf B_MIREQUESTRAMWRITEDATA139 (MIREQUESTRAMWRITEDATA[139], MIREQUESTRAMWRITEDATA_OUT[139]);
  buf B_MIREQUESTRAMWRITEDATA14 (MIREQUESTRAMWRITEDATA[14], MIREQUESTRAMWRITEDATA_OUT[14]);
  buf B_MIREQUESTRAMWRITEDATA140 (MIREQUESTRAMWRITEDATA[140], MIREQUESTRAMWRITEDATA_OUT[140]);
  buf B_MIREQUESTRAMWRITEDATA141 (MIREQUESTRAMWRITEDATA[141], MIREQUESTRAMWRITEDATA_OUT[141]);
  buf B_MIREQUESTRAMWRITEDATA142 (MIREQUESTRAMWRITEDATA[142], MIREQUESTRAMWRITEDATA_OUT[142]);
  buf B_MIREQUESTRAMWRITEDATA143 (MIREQUESTRAMWRITEDATA[143], MIREQUESTRAMWRITEDATA_OUT[143]);
  buf B_MIREQUESTRAMWRITEDATA15 (MIREQUESTRAMWRITEDATA[15], MIREQUESTRAMWRITEDATA_OUT[15]);
  buf B_MIREQUESTRAMWRITEDATA16 (MIREQUESTRAMWRITEDATA[16], MIREQUESTRAMWRITEDATA_OUT[16]);
  buf B_MIREQUESTRAMWRITEDATA17 (MIREQUESTRAMWRITEDATA[17], MIREQUESTRAMWRITEDATA_OUT[17]);
  buf B_MIREQUESTRAMWRITEDATA18 (MIREQUESTRAMWRITEDATA[18], MIREQUESTRAMWRITEDATA_OUT[18]);
  buf B_MIREQUESTRAMWRITEDATA19 (MIREQUESTRAMWRITEDATA[19], MIREQUESTRAMWRITEDATA_OUT[19]);
  buf B_MIREQUESTRAMWRITEDATA2 (MIREQUESTRAMWRITEDATA[2], MIREQUESTRAMWRITEDATA_OUT[2]);
  buf B_MIREQUESTRAMWRITEDATA20 (MIREQUESTRAMWRITEDATA[20], MIREQUESTRAMWRITEDATA_OUT[20]);
  buf B_MIREQUESTRAMWRITEDATA21 (MIREQUESTRAMWRITEDATA[21], MIREQUESTRAMWRITEDATA_OUT[21]);
  buf B_MIREQUESTRAMWRITEDATA22 (MIREQUESTRAMWRITEDATA[22], MIREQUESTRAMWRITEDATA_OUT[22]);
  buf B_MIREQUESTRAMWRITEDATA23 (MIREQUESTRAMWRITEDATA[23], MIREQUESTRAMWRITEDATA_OUT[23]);
  buf B_MIREQUESTRAMWRITEDATA24 (MIREQUESTRAMWRITEDATA[24], MIREQUESTRAMWRITEDATA_OUT[24]);
  buf B_MIREQUESTRAMWRITEDATA25 (MIREQUESTRAMWRITEDATA[25], MIREQUESTRAMWRITEDATA_OUT[25]);
  buf B_MIREQUESTRAMWRITEDATA26 (MIREQUESTRAMWRITEDATA[26], MIREQUESTRAMWRITEDATA_OUT[26]);
  buf B_MIREQUESTRAMWRITEDATA27 (MIREQUESTRAMWRITEDATA[27], MIREQUESTRAMWRITEDATA_OUT[27]);
  buf B_MIREQUESTRAMWRITEDATA28 (MIREQUESTRAMWRITEDATA[28], MIREQUESTRAMWRITEDATA_OUT[28]);
  buf B_MIREQUESTRAMWRITEDATA29 (MIREQUESTRAMWRITEDATA[29], MIREQUESTRAMWRITEDATA_OUT[29]);
  buf B_MIREQUESTRAMWRITEDATA3 (MIREQUESTRAMWRITEDATA[3], MIREQUESTRAMWRITEDATA_OUT[3]);
  buf B_MIREQUESTRAMWRITEDATA30 (MIREQUESTRAMWRITEDATA[30], MIREQUESTRAMWRITEDATA_OUT[30]);
  buf B_MIREQUESTRAMWRITEDATA31 (MIREQUESTRAMWRITEDATA[31], MIREQUESTRAMWRITEDATA_OUT[31]);
  buf B_MIREQUESTRAMWRITEDATA32 (MIREQUESTRAMWRITEDATA[32], MIREQUESTRAMWRITEDATA_OUT[32]);
  buf B_MIREQUESTRAMWRITEDATA33 (MIREQUESTRAMWRITEDATA[33], MIREQUESTRAMWRITEDATA_OUT[33]);
  buf B_MIREQUESTRAMWRITEDATA34 (MIREQUESTRAMWRITEDATA[34], MIREQUESTRAMWRITEDATA_OUT[34]);
  buf B_MIREQUESTRAMWRITEDATA35 (MIREQUESTRAMWRITEDATA[35], MIREQUESTRAMWRITEDATA_OUT[35]);
  buf B_MIREQUESTRAMWRITEDATA36 (MIREQUESTRAMWRITEDATA[36], MIREQUESTRAMWRITEDATA_OUT[36]);
  buf B_MIREQUESTRAMWRITEDATA37 (MIREQUESTRAMWRITEDATA[37], MIREQUESTRAMWRITEDATA_OUT[37]);
  buf B_MIREQUESTRAMWRITEDATA38 (MIREQUESTRAMWRITEDATA[38], MIREQUESTRAMWRITEDATA_OUT[38]);
  buf B_MIREQUESTRAMWRITEDATA39 (MIREQUESTRAMWRITEDATA[39], MIREQUESTRAMWRITEDATA_OUT[39]);
  buf B_MIREQUESTRAMWRITEDATA4 (MIREQUESTRAMWRITEDATA[4], MIREQUESTRAMWRITEDATA_OUT[4]);
  buf B_MIREQUESTRAMWRITEDATA40 (MIREQUESTRAMWRITEDATA[40], MIREQUESTRAMWRITEDATA_OUT[40]);
  buf B_MIREQUESTRAMWRITEDATA41 (MIREQUESTRAMWRITEDATA[41], MIREQUESTRAMWRITEDATA_OUT[41]);
  buf B_MIREQUESTRAMWRITEDATA42 (MIREQUESTRAMWRITEDATA[42], MIREQUESTRAMWRITEDATA_OUT[42]);
  buf B_MIREQUESTRAMWRITEDATA43 (MIREQUESTRAMWRITEDATA[43], MIREQUESTRAMWRITEDATA_OUT[43]);
  buf B_MIREQUESTRAMWRITEDATA44 (MIREQUESTRAMWRITEDATA[44], MIREQUESTRAMWRITEDATA_OUT[44]);
  buf B_MIREQUESTRAMWRITEDATA45 (MIREQUESTRAMWRITEDATA[45], MIREQUESTRAMWRITEDATA_OUT[45]);
  buf B_MIREQUESTRAMWRITEDATA46 (MIREQUESTRAMWRITEDATA[46], MIREQUESTRAMWRITEDATA_OUT[46]);
  buf B_MIREQUESTRAMWRITEDATA47 (MIREQUESTRAMWRITEDATA[47], MIREQUESTRAMWRITEDATA_OUT[47]);
  buf B_MIREQUESTRAMWRITEDATA48 (MIREQUESTRAMWRITEDATA[48], MIREQUESTRAMWRITEDATA_OUT[48]);
  buf B_MIREQUESTRAMWRITEDATA49 (MIREQUESTRAMWRITEDATA[49], MIREQUESTRAMWRITEDATA_OUT[49]);
  buf B_MIREQUESTRAMWRITEDATA5 (MIREQUESTRAMWRITEDATA[5], MIREQUESTRAMWRITEDATA_OUT[5]);
  buf B_MIREQUESTRAMWRITEDATA50 (MIREQUESTRAMWRITEDATA[50], MIREQUESTRAMWRITEDATA_OUT[50]);
  buf B_MIREQUESTRAMWRITEDATA51 (MIREQUESTRAMWRITEDATA[51], MIREQUESTRAMWRITEDATA_OUT[51]);
  buf B_MIREQUESTRAMWRITEDATA52 (MIREQUESTRAMWRITEDATA[52], MIREQUESTRAMWRITEDATA_OUT[52]);
  buf B_MIREQUESTRAMWRITEDATA53 (MIREQUESTRAMWRITEDATA[53], MIREQUESTRAMWRITEDATA_OUT[53]);
  buf B_MIREQUESTRAMWRITEDATA54 (MIREQUESTRAMWRITEDATA[54], MIREQUESTRAMWRITEDATA_OUT[54]);
  buf B_MIREQUESTRAMWRITEDATA55 (MIREQUESTRAMWRITEDATA[55], MIREQUESTRAMWRITEDATA_OUT[55]);
  buf B_MIREQUESTRAMWRITEDATA56 (MIREQUESTRAMWRITEDATA[56], MIREQUESTRAMWRITEDATA_OUT[56]);
  buf B_MIREQUESTRAMWRITEDATA57 (MIREQUESTRAMWRITEDATA[57], MIREQUESTRAMWRITEDATA_OUT[57]);
  buf B_MIREQUESTRAMWRITEDATA58 (MIREQUESTRAMWRITEDATA[58], MIREQUESTRAMWRITEDATA_OUT[58]);
  buf B_MIREQUESTRAMWRITEDATA59 (MIREQUESTRAMWRITEDATA[59], MIREQUESTRAMWRITEDATA_OUT[59]);
  buf B_MIREQUESTRAMWRITEDATA6 (MIREQUESTRAMWRITEDATA[6], MIREQUESTRAMWRITEDATA_OUT[6]);
  buf B_MIREQUESTRAMWRITEDATA60 (MIREQUESTRAMWRITEDATA[60], MIREQUESTRAMWRITEDATA_OUT[60]);
  buf B_MIREQUESTRAMWRITEDATA61 (MIREQUESTRAMWRITEDATA[61], MIREQUESTRAMWRITEDATA_OUT[61]);
  buf B_MIREQUESTRAMWRITEDATA62 (MIREQUESTRAMWRITEDATA[62], MIREQUESTRAMWRITEDATA_OUT[62]);
  buf B_MIREQUESTRAMWRITEDATA63 (MIREQUESTRAMWRITEDATA[63], MIREQUESTRAMWRITEDATA_OUT[63]);
  buf B_MIREQUESTRAMWRITEDATA64 (MIREQUESTRAMWRITEDATA[64], MIREQUESTRAMWRITEDATA_OUT[64]);
  buf B_MIREQUESTRAMWRITEDATA65 (MIREQUESTRAMWRITEDATA[65], MIREQUESTRAMWRITEDATA_OUT[65]);
  buf B_MIREQUESTRAMWRITEDATA66 (MIREQUESTRAMWRITEDATA[66], MIREQUESTRAMWRITEDATA_OUT[66]);
  buf B_MIREQUESTRAMWRITEDATA67 (MIREQUESTRAMWRITEDATA[67], MIREQUESTRAMWRITEDATA_OUT[67]);
  buf B_MIREQUESTRAMWRITEDATA68 (MIREQUESTRAMWRITEDATA[68], MIREQUESTRAMWRITEDATA_OUT[68]);
  buf B_MIREQUESTRAMWRITEDATA69 (MIREQUESTRAMWRITEDATA[69], MIREQUESTRAMWRITEDATA_OUT[69]);
  buf B_MIREQUESTRAMWRITEDATA7 (MIREQUESTRAMWRITEDATA[7], MIREQUESTRAMWRITEDATA_OUT[7]);
  buf B_MIREQUESTRAMWRITEDATA70 (MIREQUESTRAMWRITEDATA[70], MIREQUESTRAMWRITEDATA_OUT[70]);
  buf B_MIREQUESTRAMWRITEDATA71 (MIREQUESTRAMWRITEDATA[71], MIREQUESTRAMWRITEDATA_OUT[71]);
  buf B_MIREQUESTRAMWRITEDATA72 (MIREQUESTRAMWRITEDATA[72], MIREQUESTRAMWRITEDATA_OUT[72]);
  buf B_MIREQUESTRAMWRITEDATA73 (MIREQUESTRAMWRITEDATA[73], MIREQUESTRAMWRITEDATA_OUT[73]);
  buf B_MIREQUESTRAMWRITEDATA74 (MIREQUESTRAMWRITEDATA[74], MIREQUESTRAMWRITEDATA_OUT[74]);
  buf B_MIREQUESTRAMWRITEDATA75 (MIREQUESTRAMWRITEDATA[75], MIREQUESTRAMWRITEDATA_OUT[75]);
  buf B_MIREQUESTRAMWRITEDATA76 (MIREQUESTRAMWRITEDATA[76], MIREQUESTRAMWRITEDATA_OUT[76]);
  buf B_MIREQUESTRAMWRITEDATA77 (MIREQUESTRAMWRITEDATA[77], MIREQUESTRAMWRITEDATA_OUT[77]);
  buf B_MIREQUESTRAMWRITEDATA78 (MIREQUESTRAMWRITEDATA[78], MIREQUESTRAMWRITEDATA_OUT[78]);
  buf B_MIREQUESTRAMWRITEDATA79 (MIREQUESTRAMWRITEDATA[79], MIREQUESTRAMWRITEDATA_OUT[79]);
  buf B_MIREQUESTRAMWRITEDATA8 (MIREQUESTRAMWRITEDATA[8], MIREQUESTRAMWRITEDATA_OUT[8]);
  buf B_MIREQUESTRAMWRITEDATA80 (MIREQUESTRAMWRITEDATA[80], MIREQUESTRAMWRITEDATA_OUT[80]);
  buf B_MIREQUESTRAMWRITEDATA81 (MIREQUESTRAMWRITEDATA[81], MIREQUESTRAMWRITEDATA_OUT[81]);
  buf B_MIREQUESTRAMWRITEDATA82 (MIREQUESTRAMWRITEDATA[82], MIREQUESTRAMWRITEDATA_OUT[82]);
  buf B_MIREQUESTRAMWRITEDATA83 (MIREQUESTRAMWRITEDATA[83], MIREQUESTRAMWRITEDATA_OUT[83]);
  buf B_MIREQUESTRAMWRITEDATA84 (MIREQUESTRAMWRITEDATA[84], MIREQUESTRAMWRITEDATA_OUT[84]);
  buf B_MIREQUESTRAMWRITEDATA85 (MIREQUESTRAMWRITEDATA[85], MIREQUESTRAMWRITEDATA_OUT[85]);
  buf B_MIREQUESTRAMWRITEDATA86 (MIREQUESTRAMWRITEDATA[86], MIREQUESTRAMWRITEDATA_OUT[86]);
  buf B_MIREQUESTRAMWRITEDATA87 (MIREQUESTRAMWRITEDATA[87], MIREQUESTRAMWRITEDATA_OUT[87]);
  buf B_MIREQUESTRAMWRITEDATA88 (MIREQUESTRAMWRITEDATA[88], MIREQUESTRAMWRITEDATA_OUT[88]);
  buf B_MIREQUESTRAMWRITEDATA89 (MIREQUESTRAMWRITEDATA[89], MIREQUESTRAMWRITEDATA_OUT[89]);
  buf B_MIREQUESTRAMWRITEDATA9 (MIREQUESTRAMWRITEDATA[9], MIREQUESTRAMWRITEDATA_OUT[9]);
  buf B_MIREQUESTRAMWRITEDATA90 (MIREQUESTRAMWRITEDATA[90], MIREQUESTRAMWRITEDATA_OUT[90]);
  buf B_MIREQUESTRAMWRITEDATA91 (MIREQUESTRAMWRITEDATA[91], MIREQUESTRAMWRITEDATA_OUT[91]);
  buf B_MIREQUESTRAMWRITEDATA92 (MIREQUESTRAMWRITEDATA[92], MIREQUESTRAMWRITEDATA_OUT[92]);
  buf B_MIREQUESTRAMWRITEDATA93 (MIREQUESTRAMWRITEDATA[93], MIREQUESTRAMWRITEDATA_OUT[93]);
  buf B_MIREQUESTRAMWRITEDATA94 (MIREQUESTRAMWRITEDATA[94], MIREQUESTRAMWRITEDATA_OUT[94]);
  buf B_MIREQUESTRAMWRITEDATA95 (MIREQUESTRAMWRITEDATA[95], MIREQUESTRAMWRITEDATA_OUT[95]);
  buf B_MIREQUESTRAMWRITEDATA96 (MIREQUESTRAMWRITEDATA[96], MIREQUESTRAMWRITEDATA_OUT[96]);
  buf B_MIREQUESTRAMWRITEDATA97 (MIREQUESTRAMWRITEDATA[97], MIREQUESTRAMWRITEDATA_OUT[97]);
  buf B_MIREQUESTRAMWRITEDATA98 (MIREQUESTRAMWRITEDATA[98], MIREQUESTRAMWRITEDATA_OUT[98]);
  buf B_MIREQUESTRAMWRITEDATA99 (MIREQUESTRAMWRITEDATA[99], MIREQUESTRAMWRITEDATA_OUT[99]);
  buf B_MIREQUESTRAMWRITEENABLE0 (MIREQUESTRAMWRITEENABLE[0], MIREQUESTRAMWRITEENABLE_OUT[0]);
  buf B_MIREQUESTRAMWRITEENABLE1 (MIREQUESTRAMWRITEENABLE[1], MIREQUESTRAMWRITEENABLE_OUT[1]);
  buf B_MIREQUESTRAMWRITEENABLE2 (MIREQUESTRAMWRITEENABLE[2], MIREQUESTRAMWRITEENABLE_OUT[2]);
  buf B_MIREQUESTRAMWRITEENABLE3 (MIREQUESTRAMWRITEENABLE[3], MIREQUESTRAMWRITEENABLE_OUT[3]);
  buf B_PCIECQNPREQCOUNT0 (PCIECQNPREQCOUNT[0], PCIECQNPREQCOUNT_OUT[0]);
  buf B_PCIECQNPREQCOUNT1 (PCIECQNPREQCOUNT[1], PCIECQNPREQCOUNT_OUT[1]);
  buf B_PCIECQNPREQCOUNT2 (PCIECQNPREQCOUNT[2], PCIECQNPREQCOUNT_OUT[2]);
  buf B_PCIECQNPREQCOUNT3 (PCIECQNPREQCOUNT[3], PCIECQNPREQCOUNT_OUT[3]);
  buf B_PCIECQNPREQCOUNT4 (PCIECQNPREQCOUNT[4], PCIECQNPREQCOUNT_OUT[4]);
  buf B_PCIECQNPREQCOUNT5 (PCIECQNPREQCOUNT[5], PCIECQNPREQCOUNT_OUT[5]);
  buf B_PCIERQSEQNUM0 (PCIERQSEQNUM[0], PCIERQSEQNUM_OUT[0]);
  buf B_PCIERQSEQNUM1 (PCIERQSEQNUM[1], PCIERQSEQNUM_OUT[1]);
  buf B_PCIERQSEQNUM2 (PCIERQSEQNUM[2], PCIERQSEQNUM_OUT[2]);
  buf B_PCIERQSEQNUM3 (PCIERQSEQNUM[3], PCIERQSEQNUM_OUT[3]);
  buf B_PCIERQSEQNUMVLD (PCIERQSEQNUMVLD, PCIERQSEQNUMVLD_OUT);
  buf B_PCIERQTAG0 (PCIERQTAG[0], PCIERQTAG_OUT[0]);
  buf B_PCIERQTAG1 (PCIERQTAG[1], PCIERQTAG_OUT[1]);
  buf B_PCIERQTAG2 (PCIERQTAG[2], PCIERQTAG_OUT[2]);
  buf B_PCIERQTAG3 (PCIERQTAG[3], PCIERQTAG_OUT[3]);
  buf B_PCIERQTAG4 (PCIERQTAG[4], PCIERQTAG_OUT[4]);
  buf B_PCIERQTAG5 (PCIERQTAG[5], PCIERQTAG_OUT[5]);
  buf B_PCIERQTAGAV0 (PCIERQTAGAV[0], PCIERQTAGAV_OUT[0]);
  buf B_PCIERQTAGAV1 (PCIERQTAGAV[1], PCIERQTAGAV_OUT[1]);
  buf B_PCIERQTAGVLD (PCIERQTAGVLD, PCIERQTAGVLD_OUT);
  buf B_PCIETFCNPDAV0 (PCIETFCNPDAV[0], PCIETFCNPDAV_OUT[0]);
  buf B_PCIETFCNPDAV1 (PCIETFCNPDAV[1], PCIETFCNPDAV_OUT[1]);
  buf B_PCIETFCNPHAV0 (PCIETFCNPHAV[0], PCIETFCNPHAV_OUT[0]);
  buf B_PCIETFCNPHAV1 (PCIETFCNPHAV[1], PCIETFCNPHAV_OUT[1]);
  buf B_PIPERX0EQCONTROL0 (PIPERX0EQCONTROL[0], PIPERX0EQCONTROL_OUT[0]);
  buf B_PIPERX0EQCONTROL1 (PIPERX0EQCONTROL[1], PIPERX0EQCONTROL_OUT[1]);
  buf B_PIPERX0EQLPLFFS0 (PIPERX0EQLPLFFS[0], PIPERX0EQLPLFFS_OUT[0]);
  buf B_PIPERX0EQLPLFFS1 (PIPERX0EQLPLFFS[1], PIPERX0EQLPLFFS_OUT[1]);
  buf B_PIPERX0EQLPLFFS2 (PIPERX0EQLPLFFS[2], PIPERX0EQLPLFFS_OUT[2]);
  buf B_PIPERX0EQLPLFFS3 (PIPERX0EQLPLFFS[3], PIPERX0EQLPLFFS_OUT[3]);
  buf B_PIPERX0EQLPLFFS4 (PIPERX0EQLPLFFS[4], PIPERX0EQLPLFFS_OUT[4]);
  buf B_PIPERX0EQLPLFFS5 (PIPERX0EQLPLFFS[5], PIPERX0EQLPLFFS_OUT[5]);
  buf B_PIPERX0EQLPTXPRESET0 (PIPERX0EQLPTXPRESET[0], PIPERX0EQLPTXPRESET_OUT[0]);
  buf B_PIPERX0EQLPTXPRESET1 (PIPERX0EQLPTXPRESET[1], PIPERX0EQLPTXPRESET_OUT[1]);
  buf B_PIPERX0EQLPTXPRESET2 (PIPERX0EQLPTXPRESET[2], PIPERX0EQLPTXPRESET_OUT[2]);
  buf B_PIPERX0EQLPTXPRESET3 (PIPERX0EQLPTXPRESET[3], PIPERX0EQLPTXPRESET_OUT[3]);
  buf B_PIPERX0EQPRESET0 (PIPERX0EQPRESET[0], PIPERX0EQPRESET_OUT[0]);
  buf B_PIPERX0EQPRESET1 (PIPERX0EQPRESET[1], PIPERX0EQPRESET_OUT[1]);
  buf B_PIPERX0EQPRESET2 (PIPERX0EQPRESET[2], PIPERX0EQPRESET_OUT[2]);
  buf B_PIPERX0POLARITY (PIPERX0POLARITY, PIPERX0POLARITY_OUT);
  buf B_PIPERX1EQCONTROL0 (PIPERX1EQCONTROL[0], PIPERX1EQCONTROL_OUT[0]);
  buf B_PIPERX1EQCONTROL1 (PIPERX1EQCONTROL[1], PIPERX1EQCONTROL_OUT[1]);
  buf B_PIPERX1EQLPLFFS0 (PIPERX1EQLPLFFS[0], PIPERX1EQLPLFFS_OUT[0]);
  buf B_PIPERX1EQLPLFFS1 (PIPERX1EQLPLFFS[1], PIPERX1EQLPLFFS_OUT[1]);
  buf B_PIPERX1EQLPLFFS2 (PIPERX1EQLPLFFS[2], PIPERX1EQLPLFFS_OUT[2]);
  buf B_PIPERX1EQLPLFFS3 (PIPERX1EQLPLFFS[3], PIPERX1EQLPLFFS_OUT[3]);
  buf B_PIPERX1EQLPLFFS4 (PIPERX1EQLPLFFS[4], PIPERX1EQLPLFFS_OUT[4]);
  buf B_PIPERX1EQLPLFFS5 (PIPERX1EQLPLFFS[5], PIPERX1EQLPLFFS_OUT[5]);
  buf B_PIPERX1EQLPTXPRESET0 (PIPERX1EQLPTXPRESET[0], PIPERX1EQLPTXPRESET_OUT[0]);
  buf B_PIPERX1EQLPTXPRESET1 (PIPERX1EQLPTXPRESET[1], PIPERX1EQLPTXPRESET_OUT[1]);
  buf B_PIPERX1EQLPTXPRESET2 (PIPERX1EQLPTXPRESET[2], PIPERX1EQLPTXPRESET_OUT[2]);
  buf B_PIPERX1EQLPTXPRESET3 (PIPERX1EQLPTXPRESET[3], PIPERX1EQLPTXPRESET_OUT[3]);
  buf B_PIPERX1EQPRESET0 (PIPERX1EQPRESET[0], PIPERX1EQPRESET_OUT[0]);
  buf B_PIPERX1EQPRESET1 (PIPERX1EQPRESET[1], PIPERX1EQPRESET_OUT[1]);
  buf B_PIPERX1EQPRESET2 (PIPERX1EQPRESET[2], PIPERX1EQPRESET_OUT[2]);
  buf B_PIPERX1POLARITY (PIPERX1POLARITY, PIPERX1POLARITY_OUT);
  buf B_PIPERX2EQCONTROL0 (PIPERX2EQCONTROL[0], PIPERX2EQCONTROL_OUT[0]);
  buf B_PIPERX2EQCONTROL1 (PIPERX2EQCONTROL[1], PIPERX2EQCONTROL_OUT[1]);
  buf B_PIPERX2EQLPLFFS0 (PIPERX2EQLPLFFS[0], PIPERX2EQLPLFFS_OUT[0]);
  buf B_PIPERX2EQLPLFFS1 (PIPERX2EQLPLFFS[1], PIPERX2EQLPLFFS_OUT[1]);
  buf B_PIPERX2EQLPLFFS2 (PIPERX2EQLPLFFS[2], PIPERX2EQLPLFFS_OUT[2]);
  buf B_PIPERX2EQLPLFFS3 (PIPERX2EQLPLFFS[3], PIPERX2EQLPLFFS_OUT[3]);
  buf B_PIPERX2EQLPLFFS4 (PIPERX2EQLPLFFS[4], PIPERX2EQLPLFFS_OUT[4]);
  buf B_PIPERX2EQLPLFFS5 (PIPERX2EQLPLFFS[5], PIPERX2EQLPLFFS_OUT[5]);
  buf B_PIPERX2EQLPTXPRESET0 (PIPERX2EQLPTXPRESET[0], PIPERX2EQLPTXPRESET_OUT[0]);
  buf B_PIPERX2EQLPTXPRESET1 (PIPERX2EQLPTXPRESET[1], PIPERX2EQLPTXPRESET_OUT[1]);
  buf B_PIPERX2EQLPTXPRESET2 (PIPERX2EQLPTXPRESET[2], PIPERX2EQLPTXPRESET_OUT[2]);
  buf B_PIPERX2EQLPTXPRESET3 (PIPERX2EQLPTXPRESET[3], PIPERX2EQLPTXPRESET_OUT[3]);
  buf B_PIPERX2EQPRESET0 (PIPERX2EQPRESET[0], PIPERX2EQPRESET_OUT[0]);
  buf B_PIPERX2EQPRESET1 (PIPERX2EQPRESET[1], PIPERX2EQPRESET_OUT[1]);
  buf B_PIPERX2EQPRESET2 (PIPERX2EQPRESET[2], PIPERX2EQPRESET_OUT[2]);
  buf B_PIPERX2POLARITY (PIPERX2POLARITY, PIPERX2POLARITY_OUT);
  buf B_PIPERX3EQCONTROL0 (PIPERX3EQCONTROL[0], PIPERX3EQCONTROL_OUT[0]);
  buf B_PIPERX3EQCONTROL1 (PIPERX3EQCONTROL[1], PIPERX3EQCONTROL_OUT[1]);
  buf B_PIPERX3EQLPLFFS0 (PIPERX3EQLPLFFS[0], PIPERX3EQLPLFFS_OUT[0]);
  buf B_PIPERX3EQLPLFFS1 (PIPERX3EQLPLFFS[1], PIPERX3EQLPLFFS_OUT[1]);
  buf B_PIPERX3EQLPLFFS2 (PIPERX3EQLPLFFS[2], PIPERX3EQLPLFFS_OUT[2]);
  buf B_PIPERX3EQLPLFFS3 (PIPERX3EQLPLFFS[3], PIPERX3EQLPLFFS_OUT[3]);
  buf B_PIPERX3EQLPLFFS4 (PIPERX3EQLPLFFS[4], PIPERX3EQLPLFFS_OUT[4]);
  buf B_PIPERX3EQLPLFFS5 (PIPERX3EQLPLFFS[5], PIPERX3EQLPLFFS_OUT[5]);
  buf B_PIPERX3EQLPTXPRESET0 (PIPERX3EQLPTXPRESET[0], PIPERX3EQLPTXPRESET_OUT[0]);
  buf B_PIPERX3EQLPTXPRESET1 (PIPERX3EQLPTXPRESET[1], PIPERX3EQLPTXPRESET_OUT[1]);
  buf B_PIPERX3EQLPTXPRESET2 (PIPERX3EQLPTXPRESET[2], PIPERX3EQLPTXPRESET_OUT[2]);
  buf B_PIPERX3EQLPTXPRESET3 (PIPERX3EQLPTXPRESET[3], PIPERX3EQLPTXPRESET_OUT[3]);
  buf B_PIPERX3EQPRESET0 (PIPERX3EQPRESET[0], PIPERX3EQPRESET_OUT[0]);
  buf B_PIPERX3EQPRESET1 (PIPERX3EQPRESET[1], PIPERX3EQPRESET_OUT[1]);
  buf B_PIPERX3EQPRESET2 (PIPERX3EQPRESET[2], PIPERX3EQPRESET_OUT[2]);
  buf B_PIPERX3POLARITY (PIPERX3POLARITY, PIPERX3POLARITY_OUT);
  buf B_PIPERX4EQCONTROL0 (PIPERX4EQCONTROL[0], PIPERX4EQCONTROL_OUT[0]);
  buf B_PIPERX4EQCONTROL1 (PIPERX4EQCONTROL[1], PIPERX4EQCONTROL_OUT[1]);
  buf B_PIPERX4EQLPLFFS0 (PIPERX4EQLPLFFS[0], PIPERX4EQLPLFFS_OUT[0]);
  buf B_PIPERX4EQLPLFFS1 (PIPERX4EQLPLFFS[1], PIPERX4EQLPLFFS_OUT[1]);
  buf B_PIPERX4EQLPLFFS2 (PIPERX4EQLPLFFS[2], PIPERX4EQLPLFFS_OUT[2]);
  buf B_PIPERX4EQLPLFFS3 (PIPERX4EQLPLFFS[3], PIPERX4EQLPLFFS_OUT[3]);
  buf B_PIPERX4EQLPLFFS4 (PIPERX4EQLPLFFS[4], PIPERX4EQLPLFFS_OUT[4]);
  buf B_PIPERX4EQLPLFFS5 (PIPERX4EQLPLFFS[5], PIPERX4EQLPLFFS_OUT[5]);
  buf B_PIPERX4EQLPTXPRESET0 (PIPERX4EQLPTXPRESET[0], PIPERX4EQLPTXPRESET_OUT[0]);
  buf B_PIPERX4EQLPTXPRESET1 (PIPERX4EQLPTXPRESET[1], PIPERX4EQLPTXPRESET_OUT[1]);
  buf B_PIPERX4EQLPTXPRESET2 (PIPERX4EQLPTXPRESET[2], PIPERX4EQLPTXPRESET_OUT[2]);
  buf B_PIPERX4EQLPTXPRESET3 (PIPERX4EQLPTXPRESET[3], PIPERX4EQLPTXPRESET_OUT[3]);
  buf B_PIPERX4EQPRESET0 (PIPERX4EQPRESET[0], PIPERX4EQPRESET_OUT[0]);
  buf B_PIPERX4EQPRESET1 (PIPERX4EQPRESET[1], PIPERX4EQPRESET_OUT[1]);
  buf B_PIPERX4EQPRESET2 (PIPERX4EQPRESET[2], PIPERX4EQPRESET_OUT[2]);
  buf B_PIPERX4POLARITY (PIPERX4POLARITY, PIPERX4POLARITY_OUT);
  buf B_PIPERX5EQCONTROL0 (PIPERX5EQCONTROL[0], PIPERX5EQCONTROL_OUT[0]);
  buf B_PIPERX5EQCONTROL1 (PIPERX5EQCONTROL[1], PIPERX5EQCONTROL_OUT[1]);
  buf B_PIPERX5EQLPLFFS0 (PIPERX5EQLPLFFS[0], PIPERX5EQLPLFFS_OUT[0]);
  buf B_PIPERX5EQLPLFFS1 (PIPERX5EQLPLFFS[1], PIPERX5EQLPLFFS_OUT[1]);
  buf B_PIPERX5EQLPLFFS2 (PIPERX5EQLPLFFS[2], PIPERX5EQLPLFFS_OUT[2]);
  buf B_PIPERX5EQLPLFFS3 (PIPERX5EQLPLFFS[3], PIPERX5EQLPLFFS_OUT[3]);
  buf B_PIPERX5EQLPLFFS4 (PIPERX5EQLPLFFS[4], PIPERX5EQLPLFFS_OUT[4]);
  buf B_PIPERX5EQLPLFFS5 (PIPERX5EQLPLFFS[5], PIPERX5EQLPLFFS_OUT[5]);
  buf B_PIPERX5EQLPTXPRESET0 (PIPERX5EQLPTXPRESET[0], PIPERX5EQLPTXPRESET_OUT[0]);
  buf B_PIPERX5EQLPTXPRESET1 (PIPERX5EQLPTXPRESET[1], PIPERX5EQLPTXPRESET_OUT[1]);
  buf B_PIPERX5EQLPTXPRESET2 (PIPERX5EQLPTXPRESET[2], PIPERX5EQLPTXPRESET_OUT[2]);
  buf B_PIPERX5EQLPTXPRESET3 (PIPERX5EQLPTXPRESET[3], PIPERX5EQLPTXPRESET_OUT[3]);
  buf B_PIPERX5EQPRESET0 (PIPERX5EQPRESET[0], PIPERX5EQPRESET_OUT[0]);
  buf B_PIPERX5EQPRESET1 (PIPERX5EQPRESET[1], PIPERX5EQPRESET_OUT[1]);
  buf B_PIPERX5EQPRESET2 (PIPERX5EQPRESET[2], PIPERX5EQPRESET_OUT[2]);
  buf B_PIPERX5POLARITY (PIPERX5POLARITY, PIPERX5POLARITY_OUT);
  buf B_PIPERX6EQCONTROL0 (PIPERX6EQCONTROL[0], PIPERX6EQCONTROL_OUT[0]);
  buf B_PIPERX6EQCONTROL1 (PIPERX6EQCONTROL[1], PIPERX6EQCONTROL_OUT[1]);
  buf B_PIPERX6EQLPLFFS0 (PIPERX6EQLPLFFS[0], PIPERX6EQLPLFFS_OUT[0]);
  buf B_PIPERX6EQLPLFFS1 (PIPERX6EQLPLFFS[1], PIPERX6EQLPLFFS_OUT[1]);
  buf B_PIPERX6EQLPLFFS2 (PIPERX6EQLPLFFS[2], PIPERX6EQLPLFFS_OUT[2]);
  buf B_PIPERX6EQLPLFFS3 (PIPERX6EQLPLFFS[3], PIPERX6EQLPLFFS_OUT[3]);
  buf B_PIPERX6EQLPLFFS4 (PIPERX6EQLPLFFS[4], PIPERX6EQLPLFFS_OUT[4]);
  buf B_PIPERX6EQLPLFFS5 (PIPERX6EQLPLFFS[5], PIPERX6EQLPLFFS_OUT[5]);
  buf B_PIPERX6EQLPTXPRESET0 (PIPERX6EQLPTXPRESET[0], PIPERX6EQLPTXPRESET_OUT[0]);
  buf B_PIPERX6EQLPTXPRESET1 (PIPERX6EQLPTXPRESET[1], PIPERX6EQLPTXPRESET_OUT[1]);
  buf B_PIPERX6EQLPTXPRESET2 (PIPERX6EQLPTXPRESET[2], PIPERX6EQLPTXPRESET_OUT[2]);
  buf B_PIPERX6EQLPTXPRESET3 (PIPERX6EQLPTXPRESET[3], PIPERX6EQLPTXPRESET_OUT[3]);
  buf B_PIPERX6EQPRESET0 (PIPERX6EQPRESET[0], PIPERX6EQPRESET_OUT[0]);
  buf B_PIPERX6EQPRESET1 (PIPERX6EQPRESET[1], PIPERX6EQPRESET_OUT[1]);
  buf B_PIPERX6EQPRESET2 (PIPERX6EQPRESET[2], PIPERX6EQPRESET_OUT[2]);
  buf B_PIPERX6POLARITY (PIPERX6POLARITY, PIPERX6POLARITY_OUT);
  buf B_PIPERX7EQCONTROL0 (PIPERX7EQCONTROL[0], PIPERX7EQCONTROL_OUT[0]);
  buf B_PIPERX7EQCONTROL1 (PIPERX7EQCONTROL[1], PIPERX7EQCONTROL_OUT[1]);
  buf B_PIPERX7EQLPLFFS0 (PIPERX7EQLPLFFS[0], PIPERX7EQLPLFFS_OUT[0]);
  buf B_PIPERX7EQLPLFFS1 (PIPERX7EQLPLFFS[1], PIPERX7EQLPLFFS_OUT[1]);
  buf B_PIPERX7EQLPLFFS2 (PIPERX7EQLPLFFS[2], PIPERX7EQLPLFFS_OUT[2]);
  buf B_PIPERX7EQLPLFFS3 (PIPERX7EQLPLFFS[3], PIPERX7EQLPLFFS_OUT[3]);
  buf B_PIPERX7EQLPLFFS4 (PIPERX7EQLPLFFS[4], PIPERX7EQLPLFFS_OUT[4]);
  buf B_PIPERX7EQLPLFFS5 (PIPERX7EQLPLFFS[5], PIPERX7EQLPLFFS_OUT[5]);
  buf B_PIPERX7EQLPTXPRESET0 (PIPERX7EQLPTXPRESET[0], PIPERX7EQLPTXPRESET_OUT[0]);
  buf B_PIPERX7EQLPTXPRESET1 (PIPERX7EQLPTXPRESET[1], PIPERX7EQLPTXPRESET_OUT[1]);
  buf B_PIPERX7EQLPTXPRESET2 (PIPERX7EQLPTXPRESET[2], PIPERX7EQLPTXPRESET_OUT[2]);
  buf B_PIPERX7EQLPTXPRESET3 (PIPERX7EQLPTXPRESET[3], PIPERX7EQLPTXPRESET_OUT[3]);
  buf B_PIPERX7EQPRESET0 (PIPERX7EQPRESET[0], PIPERX7EQPRESET_OUT[0]);
  buf B_PIPERX7EQPRESET1 (PIPERX7EQPRESET[1], PIPERX7EQPRESET_OUT[1]);
  buf B_PIPERX7EQPRESET2 (PIPERX7EQPRESET[2], PIPERX7EQPRESET_OUT[2]);
  buf B_PIPERX7POLARITY (PIPERX7POLARITY, PIPERX7POLARITY_OUT);
  buf B_PIPETX0CHARISK0 (PIPETX0CHARISK[0], PIPETX0CHARISK_OUT[0]);
  buf B_PIPETX0CHARISK1 (PIPETX0CHARISK[1], PIPETX0CHARISK_OUT[1]);
  buf B_PIPETX0COMPLIANCE (PIPETX0COMPLIANCE, PIPETX0COMPLIANCE_OUT);
  buf B_PIPETX0DATA0 (PIPETX0DATA[0], PIPETX0DATA_OUT[0]);
  buf B_PIPETX0DATA1 (PIPETX0DATA[1], PIPETX0DATA_OUT[1]);
  buf B_PIPETX0DATA10 (PIPETX0DATA[10], PIPETX0DATA_OUT[10]);
  buf B_PIPETX0DATA11 (PIPETX0DATA[11], PIPETX0DATA_OUT[11]);
  buf B_PIPETX0DATA12 (PIPETX0DATA[12], PIPETX0DATA_OUT[12]);
  buf B_PIPETX0DATA13 (PIPETX0DATA[13], PIPETX0DATA_OUT[13]);
  buf B_PIPETX0DATA14 (PIPETX0DATA[14], PIPETX0DATA_OUT[14]);
  buf B_PIPETX0DATA15 (PIPETX0DATA[15], PIPETX0DATA_OUT[15]);
  buf B_PIPETX0DATA16 (PIPETX0DATA[16], PIPETX0DATA_OUT[16]);
  buf B_PIPETX0DATA17 (PIPETX0DATA[17], PIPETX0DATA_OUT[17]);
  buf B_PIPETX0DATA18 (PIPETX0DATA[18], PIPETX0DATA_OUT[18]);
  buf B_PIPETX0DATA19 (PIPETX0DATA[19], PIPETX0DATA_OUT[19]);
  buf B_PIPETX0DATA2 (PIPETX0DATA[2], PIPETX0DATA_OUT[2]);
  buf B_PIPETX0DATA20 (PIPETX0DATA[20], PIPETX0DATA_OUT[20]);
  buf B_PIPETX0DATA21 (PIPETX0DATA[21], PIPETX0DATA_OUT[21]);
  buf B_PIPETX0DATA22 (PIPETX0DATA[22], PIPETX0DATA_OUT[22]);
  buf B_PIPETX0DATA23 (PIPETX0DATA[23], PIPETX0DATA_OUT[23]);
  buf B_PIPETX0DATA24 (PIPETX0DATA[24], PIPETX0DATA_OUT[24]);
  buf B_PIPETX0DATA25 (PIPETX0DATA[25], PIPETX0DATA_OUT[25]);
  buf B_PIPETX0DATA26 (PIPETX0DATA[26], PIPETX0DATA_OUT[26]);
  buf B_PIPETX0DATA27 (PIPETX0DATA[27], PIPETX0DATA_OUT[27]);
  buf B_PIPETX0DATA28 (PIPETX0DATA[28], PIPETX0DATA_OUT[28]);
  buf B_PIPETX0DATA29 (PIPETX0DATA[29], PIPETX0DATA_OUT[29]);
  buf B_PIPETX0DATA3 (PIPETX0DATA[3], PIPETX0DATA_OUT[3]);
  buf B_PIPETX0DATA30 (PIPETX0DATA[30], PIPETX0DATA_OUT[30]);
  buf B_PIPETX0DATA31 (PIPETX0DATA[31], PIPETX0DATA_OUT[31]);
  buf B_PIPETX0DATA4 (PIPETX0DATA[4], PIPETX0DATA_OUT[4]);
  buf B_PIPETX0DATA5 (PIPETX0DATA[5], PIPETX0DATA_OUT[5]);
  buf B_PIPETX0DATA6 (PIPETX0DATA[6], PIPETX0DATA_OUT[6]);
  buf B_PIPETX0DATA7 (PIPETX0DATA[7], PIPETX0DATA_OUT[7]);
  buf B_PIPETX0DATA8 (PIPETX0DATA[8], PIPETX0DATA_OUT[8]);
  buf B_PIPETX0DATA9 (PIPETX0DATA[9], PIPETX0DATA_OUT[9]);
  buf B_PIPETX0DATAVALID (PIPETX0DATAVALID, PIPETX0DATAVALID_OUT);
  buf B_PIPETX0ELECIDLE (PIPETX0ELECIDLE, PIPETX0ELECIDLE_OUT);
  buf B_PIPETX0EQCONTROL0 (PIPETX0EQCONTROL[0], PIPETX0EQCONTROL_OUT[0]);
  buf B_PIPETX0EQCONTROL1 (PIPETX0EQCONTROL[1], PIPETX0EQCONTROL_OUT[1]);
  buf B_PIPETX0EQDEEMPH0 (PIPETX0EQDEEMPH[0], PIPETX0EQDEEMPH_OUT[0]);
  buf B_PIPETX0EQDEEMPH1 (PIPETX0EQDEEMPH[1], PIPETX0EQDEEMPH_OUT[1]);
  buf B_PIPETX0EQDEEMPH2 (PIPETX0EQDEEMPH[2], PIPETX0EQDEEMPH_OUT[2]);
  buf B_PIPETX0EQDEEMPH3 (PIPETX0EQDEEMPH[3], PIPETX0EQDEEMPH_OUT[3]);
  buf B_PIPETX0EQDEEMPH4 (PIPETX0EQDEEMPH[4], PIPETX0EQDEEMPH_OUT[4]);
  buf B_PIPETX0EQDEEMPH5 (PIPETX0EQDEEMPH[5], PIPETX0EQDEEMPH_OUT[5]);
  buf B_PIPETX0EQPRESET0 (PIPETX0EQPRESET[0], PIPETX0EQPRESET_OUT[0]);
  buf B_PIPETX0EQPRESET1 (PIPETX0EQPRESET[1], PIPETX0EQPRESET_OUT[1]);
  buf B_PIPETX0EQPRESET2 (PIPETX0EQPRESET[2], PIPETX0EQPRESET_OUT[2]);
  buf B_PIPETX0EQPRESET3 (PIPETX0EQPRESET[3], PIPETX0EQPRESET_OUT[3]);
  buf B_PIPETX0POWERDOWN0 (PIPETX0POWERDOWN[0], PIPETX0POWERDOWN_OUT[0]);
  buf B_PIPETX0POWERDOWN1 (PIPETX0POWERDOWN[1], PIPETX0POWERDOWN_OUT[1]);
  buf B_PIPETX0STARTBLOCK (PIPETX0STARTBLOCK, PIPETX0STARTBLOCK_OUT);
  buf B_PIPETX0SYNCHEADER0 (PIPETX0SYNCHEADER[0], PIPETX0SYNCHEADER_OUT[0]);
  buf B_PIPETX0SYNCHEADER1 (PIPETX0SYNCHEADER[1], PIPETX0SYNCHEADER_OUT[1]);
  buf B_PIPETX1CHARISK0 (PIPETX1CHARISK[0], PIPETX1CHARISK_OUT[0]);
  buf B_PIPETX1CHARISK1 (PIPETX1CHARISK[1], PIPETX1CHARISK_OUT[1]);
  buf B_PIPETX1COMPLIANCE (PIPETX1COMPLIANCE, PIPETX1COMPLIANCE_OUT);
  buf B_PIPETX1DATA0 (PIPETX1DATA[0], PIPETX1DATA_OUT[0]);
  buf B_PIPETX1DATA1 (PIPETX1DATA[1], PIPETX1DATA_OUT[1]);
  buf B_PIPETX1DATA10 (PIPETX1DATA[10], PIPETX1DATA_OUT[10]);
  buf B_PIPETX1DATA11 (PIPETX1DATA[11], PIPETX1DATA_OUT[11]);
  buf B_PIPETX1DATA12 (PIPETX1DATA[12], PIPETX1DATA_OUT[12]);
  buf B_PIPETX1DATA13 (PIPETX1DATA[13], PIPETX1DATA_OUT[13]);
  buf B_PIPETX1DATA14 (PIPETX1DATA[14], PIPETX1DATA_OUT[14]);
  buf B_PIPETX1DATA15 (PIPETX1DATA[15], PIPETX1DATA_OUT[15]);
  buf B_PIPETX1DATA16 (PIPETX1DATA[16], PIPETX1DATA_OUT[16]);
  buf B_PIPETX1DATA17 (PIPETX1DATA[17], PIPETX1DATA_OUT[17]);
  buf B_PIPETX1DATA18 (PIPETX1DATA[18], PIPETX1DATA_OUT[18]);
  buf B_PIPETX1DATA19 (PIPETX1DATA[19], PIPETX1DATA_OUT[19]);
  buf B_PIPETX1DATA2 (PIPETX1DATA[2], PIPETX1DATA_OUT[2]);
  buf B_PIPETX1DATA20 (PIPETX1DATA[20], PIPETX1DATA_OUT[20]);
  buf B_PIPETX1DATA21 (PIPETX1DATA[21], PIPETX1DATA_OUT[21]);
  buf B_PIPETX1DATA22 (PIPETX1DATA[22], PIPETX1DATA_OUT[22]);
  buf B_PIPETX1DATA23 (PIPETX1DATA[23], PIPETX1DATA_OUT[23]);
  buf B_PIPETX1DATA24 (PIPETX1DATA[24], PIPETX1DATA_OUT[24]);
  buf B_PIPETX1DATA25 (PIPETX1DATA[25], PIPETX1DATA_OUT[25]);
  buf B_PIPETX1DATA26 (PIPETX1DATA[26], PIPETX1DATA_OUT[26]);
  buf B_PIPETX1DATA27 (PIPETX1DATA[27], PIPETX1DATA_OUT[27]);
  buf B_PIPETX1DATA28 (PIPETX1DATA[28], PIPETX1DATA_OUT[28]);
  buf B_PIPETX1DATA29 (PIPETX1DATA[29], PIPETX1DATA_OUT[29]);
  buf B_PIPETX1DATA3 (PIPETX1DATA[3], PIPETX1DATA_OUT[3]);
  buf B_PIPETX1DATA30 (PIPETX1DATA[30], PIPETX1DATA_OUT[30]);
  buf B_PIPETX1DATA31 (PIPETX1DATA[31], PIPETX1DATA_OUT[31]);
  buf B_PIPETX1DATA4 (PIPETX1DATA[4], PIPETX1DATA_OUT[4]);
  buf B_PIPETX1DATA5 (PIPETX1DATA[5], PIPETX1DATA_OUT[5]);
  buf B_PIPETX1DATA6 (PIPETX1DATA[6], PIPETX1DATA_OUT[6]);
  buf B_PIPETX1DATA7 (PIPETX1DATA[7], PIPETX1DATA_OUT[7]);
  buf B_PIPETX1DATA8 (PIPETX1DATA[8], PIPETX1DATA_OUT[8]);
  buf B_PIPETX1DATA9 (PIPETX1DATA[9], PIPETX1DATA_OUT[9]);
  buf B_PIPETX1DATAVALID (PIPETX1DATAVALID, PIPETX1DATAVALID_OUT);
  buf B_PIPETX1ELECIDLE (PIPETX1ELECIDLE, PIPETX1ELECIDLE_OUT);
  buf B_PIPETX1EQCONTROL0 (PIPETX1EQCONTROL[0], PIPETX1EQCONTROL_OUT[0]);
  buf B_PIPETX1EQCONTROL1 (PIPETX1EQCONTROL[1], PIPETX1EQCONTROL_OUT[1]);
  buf B_PIPETX1EQDEEMPH0 (PIPETX1EQDEEMPH[0], PIPETX1EQDEEMPH_OUT[0]);
  buf B_PIPETX1EQDEEMPH1 (PIPETX1EQDEEMPH[1], PIPETX1EQDEEMPH_OUT[1]);
  buf B_PIPETX1EQDEEMPH2 (PIPETX1EQDEEMPH[2], PIPETX1EQDEEMPH_OUT[2]);
  buf B_PIPETX1EQDEEMPH3 (PIPETX1EQDEEMPH[3], PIPETX1EQDEEMPH_OUT[3]);
  buf B_PIPETX1EQDEEMPH4 (PIPETX1EQDEEMPH[4], PIPETX1EQDEEMPH_OUT[4]);
  buf B_PIPETX1EQDEEMPH5 (PIPETX1EQDEEMPH[5], PIPETX1EQDEEMPH_OUT[5]);
  buf B_PIPETX1EQPRESET0 (PIPETX1EQPRESET[0], PIPETX1EQPRESET_OUT[0]);
  buf B_PIPETX1EQPRESET1 (PIPETX1EQPRESET[1], PIPETX1EQPRESET_OUT[1]);
  buf B_PIPETX1EQPRESET2 (PIPETX1EQPRESET[2], PIPETX1EQPRESET_OUT[2]);
  buf B_PIPETX1EQPRESET3 (PIPETX1EQPRESET[3], PIPETX1EQPRESET_OUT[3]);
  buf B_PIPETX1POWERDOWN0 (PIPETX1POWERDOWN[0], PIPETX1POWERDOWN_OUT[0]);
  buf B_PIPETX1POWERDOWN1 (PIPETX1POWERDOWN[1], PIPETX1POWERDOWN_OUT[1]);
  buf B_PIPETX1STARTBLOCK (PIPETX1STARTBLOCK, PIPETX1STARTBLOCK_OUT);
  buf B_PIPETX1SYNCHEADER0 (PIPETX1SYNCHEADER[0], PIPETX1SYNCHEADER_OUT[0]);
  buf B_PIPETX1SYNCHEADER1 (PIPETX1SYNCHEADER[1], PIPETX1SYNCHEADER_OUT[1]);
  buf B_PIPETX2CHARISK0 (PIPETX2CHARISK[0], PIPETX2CHARISK_OUT[0]);
  buf B_PIPETX2CHARISK1 (PIPETX2CHARISK[1], PIPETX2CHARISK_OUT[1]);
  buf B_PIPETX2COMPLIANCE (PIPETX2COMPLIANCE, PIPETX2COMPLIANCE_OUT);
  buf B_PIPETX2DATA0 (PIPETX2DATA[0], PIPETX2DATA_OUT[0]);
  buf B_PIPETX2DATA1 (PIPETX2DATA[1], PIPETX2DATA_OUT[1]);
  buf B_PIPETX2DATA10 (PIPETX2DATA[10], PIPETX2DATA_OUT[10]);
  buf B_PIPETX2DATA11 (PIPETX2DATA[11], PIPETX2DATA_OUT[11]);
  buf B_PIPETX2DATA12 (PIPETX2DATA[12], PIPETX2DATA_OUT[12]);
  buf B_PIPETX2DATA13 (PIPETX2DATA[13], PIPETX2DATA_OUT[13]);
  buf B_PIPETX2DATA14 (PIPETX2DATA[14], PIPETX2DATA_OUT[14]);
  buf B_PIPETX2DATA15 (PIPETX2DATA[15], PIPETX2DATA_OUT[15]);
  buf B_PIPETX2DATA16 (PIPETX2DATA[16], PIPETX2DATA_OUT[16]);
  buf B_PIPETX2DATA17 (PIPETX2DATA[17], PIPETX2DATA_OUT[17]);
  buf B_PIPETX2DATA18 (PIPETX2DATA[18], PIPETX2DATA_OUT[18]);
  buf B_PIPETX2DATA19 (PIPETX2DATA[19], PIPETX2DATA_OUT[19]);
  buf B_PIPETX2DATA2 (PIPETX2DATA[2], PIPETX2DATA_OUT[2]);
  buf B_PIPETX2DATA20 (PIPETX2DATA[20], PIPETX2DATA_OUT[20]);
  buf B_PIPETX2DATA21 (PIPETX2DATA[21], PIPETX2DATA_OUT[21]);
  buf B_PIPETX2DATA22 (PIPETX2DATA[22], PIPETX2DATA_OUT[22]);
  buf B_PIPETX2DATA23 (PIPETX2DATA[23], PIPETX2DATA_OUT[23]);
  buf B_PIPETX2DATA24 (PIPETX2DATA[24], PIPETX2DATA_OUT[24]);
  buf B_PIPETX2DATA25 (PIPETX2DATA[25], PIPETX2DATA_OUT[25]);
  buf B_PIPETX2DATA26 (PIPETX2DATA[26], PIPETX2DATA_OUT[26]);
  buf B_PIPETX2DATA27 (PIPETX2DATA[27], PIPETX2DATA_OUT[27]);
  buf B_PIPETX2DATA28 (PIPETX2DATA[28], PIPETX2DATA_OUT[28]);
  buf B_PIPETX2DATA29 (PIPETX2DATA[29], PIPETX2DATA_OUT[29]);
  buf B_PIPETX2DATA3 (PIPETX2DATA[3], PIPETX2DATA_OUT[3]);
  buf B_PIPETX2DATA30 (PIPETX2DATA[30], PIPETX2DATA_OUT[30]);
  buf B_PIPETX2DATA31 (PIPETX2DATA[31], PIPETX2DATA_OUT[31]);
  buf B_PIPETX2DATA4 (PIPETX2DATA[4], PIPETX2DATA_OUT[4]);
  buf B_PIPETX2DATA5 (PIPETX2DATA[5], PIPETX2DATA_OUT[5]);
  buf B_PIPETX2DATA6 (PIPETX2DATA[6], PIPETX2DATA_OUT[6]);
  buf B_PIPETX2DATA7 (PIPETX2DATA[7], PIPETX2DATA_OUT[7]);
  buf B_PIPETX2DATA8 (PIPETX2DATA[8], PIPETX2DATA_OUT[8]);
  buf B_PIPETX2DATA9 (PIPETX2DATA[9], PIPETX2DATA_OUT[9]);
  buf B_PIPETX2DATAVALID (PIPETX2DATAVALID, PIPETX2DATAVALID_OUT);
  buf B_PIPETX2ELECIDLE (PIPETX2ELECIDLE, PIPETX2ELECIDLE_OUT);
  buf B_PIPETX2EQCONTROL0 (PIPETX2EQCONTROL[0], PIPETX2EQCONTROL_OUT[0]);
  buf B_PIPETX2EQCONTROL1 (PIPETX2EQCONTROL[1], PIPETX2EQCONTROL_OUT[1]);
  buf B_PIPETX2EQDEEMPH0 (PIPETX2EQDEEMPH[0], PIPETX2EQDEEMPH_OUT[0]);
  buf B_PIPETX2EQDEEMPH1 (PIPETX2EQDEEMPH[1], PIPETX2EQDEEMPH_OUT[1]);
  buf B_PIPETX2EQDEEMPH2 (PIPETX2EQDEEMPH[2], PIPETX2EQDEEMPH_OUT[2]);
  buf B_PIPETX2EQDEEMPH3 (PIPETX2EQDEEMPH[3], PIPETX2EQDEEMPH_OUT[3]);
  buf B_PIPETX2EQDEEMPH4 (PIPETX2EQDEEMPH[4], PIPETX2EQDEEMPH_OUT[4]);
  buf B_PIPETX2EQDEEMPH5 (PIPETX2EQDEEMPH[5], PIPETX2EQDEEMPH_OUT[5]);
  buf B_PIPETX2EQPRESET0 (PIPETX2EQPRESET[0], PIPETX2EQPRESET_OUT[0]);
  buf B_PIPETX2EQPRESET1 (PIPETX2EQPRESET[1], PIPETX2EQPRESET_OUT[1]);
  buf B_PIPETX2EQPRESET2 (PIPETX2EQPRESET[2], PIPETX2EQPRESET_OUT[2]);
  buf B_PIPETX2EQPRESET3 (PIPETX2EQPRESET[3], PIPETX2EQPRESET_OUT[3]);
  buf B_PIPETX2POWERDOWN0 (PIPETX2POWERDOWN[0], PIPETX2POWERDOWN_OUT[0]);
  buf B_PIPETX2POWERDOWN1 (PIPETX2POWERDOWN[1], PIPETX2POWERDOWN_OUT[1]);
  buf B_PIPETX2STARTBLOCK (PIPETX2STARTBLOCK, PIPETX2STARTBLOCK_OUT);
  buf B_PIPETX2SYNCHEADER0 (PIPETX2SYNCHEADER[0], PIPETX2SYNCHEADER_OUT[0]);
  buf B_PIPETX2SYNCHEADER1 (PIPETX2SYNCHEADER[1], PIPETX2SYNCHEADER_OUT[1]);
  buf B_PIPETX3CHARISK0 (PIPETX3CHARISK[0], PIPETX3CHARISK_OUT[0]);
  buf B_PIPETX3CHARISK1 (PIPETX3CHARISK[1], PIPETX3CHARISK_OUT[1]);
  buf B_PIPETX3COMPLIANCE (PIPETX3COMPLIANCE, PIPETX3COMPLIANCE_OUT);
  buf B_PIPETX3DATA0 (PIPETX3DATA[0], PIPETX3DATA_OUT[0]);
  buf B_PIPETX3DATA1 (PIPETX3DATA[1], PIPETX3DATA_OUT[1]);
  buf B_PIPETX3DATA10 (PIPETX3DATA[10], PIPETX3DATA_OUT[10]);
  buf B_PIPETX3DATA11 (PIPETX3DATA[11], PIPETX3DATA_OUT[11]);
  buf B_PIPETX3DATA12 (PIPETX3DATA[12], PIPETX3DATA_OUT[12]);
  buf B_PIPETX3DATA13 (PIPETX3DATA[13], PIPETX3DATA_OUT[13]);
  buf B_PIPETX3DATA14 (PIPETX3DATA[14], PIPETX3DATA_OUT[14]);
  buf B_PIPETX3DATA15 (PIPETX3DATA[15], PIPETX3DATA_OUT[15]);
  buf B_PIPETX3DATA16 (PIPETX3DATA[16], PIPETX3DATA_OUT[16]);
  buf B_PIPETX3DATA17 (PIPETX3DATA[17], PIPETX3DATA_OUT[17]);
  buf B_PIPETX3DATA18 (PIPETX3DATA[18], PIPETX3DATA_OUT[18]);
  buf B_PIPETX3DATA19 (PIPETX3DATA[19], PIPETX3DATA_OUT[19]);
  buf B_PIPETX3DATA2 (PIPETX3DATA[2], PIPETX3DATA_OUT[2]);
  buf B_PIPETX3DATA20 (PIPETX3DATA[20], PIPETX3DATA_OUT[20]);
  buf B_PIPETX3DATA21 (PIPETX3DATA[21], PIPETX3DATA_OUT[21]);
  buf B_PIPETX3DATA22 (PIPETX3DATA[22], PIPETX3DATA_OUT[22]);
  buf B_PIPETX3DATA23 (PIPETX3DATA[23], PIPETX3DATA_OUT[23]);
  buf B_PIPETX3DATA24 (PIPETX3DATA[24], PIPETX3DATA_OUT[24]);
  buf B_PIPETX3DATA25 (PIPETX3DATA[25], PIPETX3DATA_OUT[25]);
  buf B_PIPETX3DATA26 (PIPETX3DATA[26], PIPETX3DATA_OUT[26]);
  buf B_PIPETX3DATA27 (PIPETX3DATA[27], PIPETX3DATA_OUT[27]);
  buf B_PIPETX3DATA28 (PIPETX3DATA[28], PIPETX3DATA_OUT[28]);
  buf B_PIPETX3DATA29 (PIPETX3DATA[29], PIPETX3DATA_OUT[29]);
  buf B_PIPETX3DATA3 (PIPETX3DATA[3], PIPETX3DATA_OUT[3]);
  buf B_PIPETX3DATA30 (PIPETX3DATA[30], PIPETX3DATA_OUT[30]);
  buf B_PIPETX3DATA31 (PIPETX3DATA[31], PIPETX3DATA_OUT[31]);
  buf B_PIPETX3DATA4 (PIPETX3DATA[4], PIPETX3DATA_OUT[4]);
  buf B_PIPETX3DATA5 (PIPETX3DATA[5], PIPETX3DATA_OUT[5]);
  buf B_PIPETX3DATA6 (PIPETX3DATA[6], PIPETX3DATA_OUT[6]);
  buf B_PIPETX3DATA7 (PIPETX3DATA[7], PIPETX3DATA_OUT[7]);
  buf B_PIPETX3DATA8 (PIPETX3DATA[8], PIPETX3DATA_OUT[8]);
  buf B_PIPETX3DATA9 (PIPETX3DATA[9], PIPETX3DATA_OUT[9]);
  buf B_PIPETX3DATAVALID (PIPETX3DATAVALID, PIPETX3DATAVALID_OUT);
  buf B_PIPETX3ELECIDLE (PIPETX3ELECIDLE, PIPETX3ELECIDLE_OUT);
  buf B_PIPETX3EQCONTROL0 (PIPETX3EQCONTROL[0], PIPETX3EQCONTROL_OUT[0]);
  buf B_PIPETX3EQCONTROL1 (PIPETX3EQCONTROL[1], PIPETX3EQCONTROL_OUT[1]);
  buf B_PIPETX3EQDEEMPH0 (PIPETX3EQDEEMPH[0], PIPETX3EQDEEMPH_OUT[0]);
  buf B_PIPETX3EQDEEMPH1 (PIPETX3EQDEEMPH[1], PIPETX3EQDEEMPH_OUT[1]);
  buf B_PIPETX3EQDEEMPH2 (PIPETX3EQDEEMPH[2], PIPETX3EQDEEMPH_OUT[2]);
  buf B_PIPETX3EQDEEMPH3 (PIPETX3EQDEEMPH[3], PIPETX3EQDEEMPH_OUT[3]);
  buf B_PIPETX3EQDEEMPH4 (PIPETX3EQDEEMPH[4], PIPETX3EQDEEMPH_OUT[4]);
  buf B_PIPETX3EQDEEMPH5 (PIPETX3EQDEEMPH[5], PIPETX3EQDEEMPH_OUT[5]);
  buf B_PIPETX3EQPRESET0 (PIPETX3EQPRESET[0], PIPETX3EQPRESET_OUT[0]);
  buf B_PIPETX3EQPRESET1 (PIPETX3EQPRESET[1], PIPETX3EQPRESET_OUT[1]);
  buf B_PIPETX3EQPRESET2 (PIPETX3EQPRESET[2], PIPETX3EQPRESET_OUT[2]);
  buf B_PIPETX3EQPRESET3 (PIPETX3EQPRESET[3], PIPETX3EQPRESET_OUT[3]);
  buf B_PIPETX3POWERDOWN0 (PIPETX3POWERDOWN[0], PIPETX3POWERDOWN_OUT[0]);
  buf B_PIPETX3POWERDOWN1 (PIPETX3POWERDOWN[1], PIPETX3POWERDOWN_OUT[1]);
  buf B_PIPETX3STARTBLOCK (PIPETX3STARTBLOCK, PIPETX3STARTBLOCK_OUT);
  buf B_PIPETX3SYNCHEADER0 (PIPETX3SYNCHEADER[0], PIPETX3SYNCHEADER_OUT[0]);
  buf B_PIPETX3SYNCHEADER1 (PIPETX3SYNCHEADER[1], PIPETX3SYNCHEADER_OUT[1]);
  buf B_PIPETX4CHARISK0 (PIPETX4CHARISK[0], PIPETX4CHARISK_OUT[0]);
  buf B_PIPETX4CHARISK1 (PIPETX4CHARISK[1], PIPETX4CHARISK_OUT[1]);
  buf B_PIPETX4COMPLIANCE (PIPETX4COMPLIANCE, PIPETX4COMPLIANCE_OUT);
  buf B_PIPETX4DATA0 (PIPETX4DATA[0], PIPETX4DATA_OUT[0]);
  buf B_PIPETX4DATA1 (PIPETX4DATA[1], PIPETX4DATA_OUT[1]);
  buf B_PIPETX4DATA10 (PIPETX4DATA[10], PIPETX4DATA_OUT[10]);
  buf B_PIPETX4DATA11 (PIPETX4DATA[11], PIPETX4DATA_OUT[11]);
  buf B_PIPETX4DATA12 (PIPETX4DATA[12], PIPETX4DATA_OUT[12]);
  buf B_PIPETX4DATA13 (PIPETX4DATA[13], PIPETX4DATA_OUT[13]);
  buf B_PIPETX4DATA14 (PIPETX4DATA[14], PIPETX4DATA_OUT[14]);
  buf B_PIPETX4DATA15 (PIPETX4DATA[15], PIPETX4DATA_OUT[15]);
  buf B_PIPETX4DATA16 (PIPETX4DATA[16], PIPETX4DATA_OUT[16]);
  buf B_PIPETX4DATA17 (PIPETX4DATA[17], PIPETX4DATA_OUT[17]);
  buf B_PIPETX4DATA18 (PIPETX4DATA[18], PIPETX4DATA_OUT[18]);
  buf B_PIPETX4DATA19 (PIPETX4DATA[19], PIPETX4DATA_OUT[19]);
  buf B_PIPETX4DATA2 (PIPETX4DATA[2], PIPETX4DATA_OUT[2]);
  buf B_PIPETX4DATA20 (PIPETX4DATA[20], PIPETX4DATA_OUT[20]);
  buf B_PIPETX4DATA21 (PIPETX4DATA[21], PIPETX4DATA_OUT[21]);
  buf B_PIPETX4DATA22 (PIPETX4DATA[22], PIPETX4DATA_OUT[22]);
  buf B_PIPETX4DATA23 (PIPETX4DATA[23], PIPETX4DATA_OUT[23]);
  buf B_PIPETX4DATA24 (PIPETX4DATA[24], PIPETX4DATA_OUT[24]);
  buf B_PIPETX4DATA25 (PIPETX4DATA[25], PIPETX4DATA_OUT[25]);
  buf B_PIPETX4DATA26 (PIPETX4DATA[26], PIPETX4DATA_OUT[26]);
  buf B_PIPETX4DATA27 (PIPETX4DATA[27], PIPETX4DATA_OUT[27]);
  buf B_PIPETX4DATA28 (PIPETX4DATA[28], PIPETX4DATA_OUT[28]);
  buf B_PIPETX4DATA29 (PIPETX4DATA[29], PIPETX4DATA_OUT[29]);
  buf B_PIPETX4DATA3 (PIPETX4DATA[3], PIPETX4DATA_OUT[3]);
  buf B_PIPETX4DATA30 (PIPETX4DATA[30], PIPETX4DATA_OUT[30]);
  buf B_PIPETX4DATA31 (PIPETX4DATA[31], PIPETX4DATA_OUT[31]);
  buf B_PIPETX4DATA4 (PIPETX4DATA[4], PIPETX4DATA_OUT[4]);
  buf B_PIPETX4DATA5 (PIPETX4DATA[5], PIPETX4DATA_OUT[5]);
  buf B_PIPETX4DATA6 (PIPETX4DATA[6], PIPETX4DATA_OUT[6]);
  buf B_PIPETX4DATA7 (PIPETX4DATA[7], PIPETX4DATA_OUT[7]);
  buf B_PIPETX4DATA8 (PIPETX4DATA[8], PIPETX4DATA_OUT[8]);
  buf B_PIPETX4DATA9 (PIPETX4DATA[9], PIPETX4DATA_OUT[9]);
  buf B_PIPETX4DATAVALID (PIPETX4DATAVALID, PIPETX4DATAVALID_OUT);
  buf B_PIPETX4ELECIDLE (PIPETX4ELECIDLE, PIPETX4ELECIDLE_OUT);
  buf B_PIPETX4EQCONTROL0 (PIPETX4EQCONTROL[0], PIPETX4EQCONTROL_OUT[0]);
  buf B_PIPETX4EQCONTROL1 (PIPETX4EQCONTROL[1], PIPETX4EQCONTROL_OUT[1]);
  buf B_PIPETX4EQDEEMPH0 (PIPETX4EQDEEMPH[0], PIPETX4EQDEEMPH_OUT[0]);
  buf B_PIPETX4EQDEEMPH1 (PIPETX4EQDEEMPH[1], PIPETX4EQDEEMPH_OUT[1]);
  buf B_PIPETX4EQDEEMPH2 (PIPETX4EQDEEMPH[2], PIPETX4EQDEEMPH_OUT[2]);
  buf B_PIPETX4EQDEEMPH3 (PIPETX4EQDEEMPH[3], PIPETX4EQDEEMPH_OUT[3]);
  buf B_PIPETX4EQDEEMPH4 (PIPETX4EQDEEMPH[4], PIPETX4EQDEEMPH_OUT[4]);
  buf B_PIPETX4EQDEEMPH5 (PIPETX4EQDEEMPH[5], PIPETX4EQDEEMPH_OUT[5]);
  buf B_PIPETX4EQPRESET0 (PIPETX4EQPRESET[0], PIPETX4EQPRESET_OUT[0]);
  buf B_PIPETX4EQPRESET1 (PIPETX4EQPRESET[1], PIPETX4EQPRESET_OUT[1]);
  buf B_PIPETX4EQPRESET2 (PIPETX4EQPRESET[2], PIPETX4EQPRESET_OUT[2]);
  buf B_PIPETX4EQPRESET3 (PIPETX4EQPRESET[3], PIPETX4EQPRESET_OUT[3]);
  buf B_PIPETX4POWERDOWN0 (PIPETX4POWERDOWN[0], PIPETX4POWERDOWN_OUT[0]);
  buf B_PIPETX4POWERDOWN1 (PIPETX4POWERDOWN[1], PIPETX4POWERDOWN_OUT[1]);
  buf B_PIPETX4STARTBLOCK (PIPETX4STARTBLOCK, PIPETX4STARTBLOCK_OUT);
  buf B_PIPETX4SYNCHEADER0 (PIPETX4SYNCHEADER[0], PIPETX4SYNCHEADER_OUT[0]);
  buf B_PIPETX4SYNCHEADER1 (PIPETX4SYNCHEADER[1], PIPETX4SYNCHEADER_OUT[1]);
  buf B_PIPETX5CHARISK0 (PIPETX5CHARISK[0], PIPETX5CHARISK_OUT[0]);
  buf B_PIPETX5CHARISK1 (PIPETX5CHARISK[1], PIPETX5CHARISK_OUT[1]);
  buf B_PIPETX5COMPLIANCE (PIPETX5COMPLIANCE, PIPETX5COMPLIANCE_OUT);
  buf B_PIPETX5DATA0 (PIPETX5DATA[0], PIPETX5DATA_OUT[0]);
  buf B_PIPETX5DATA1 (PIPETX5DATA[1], PIPETX5DATA_OUT[1]);
  buf B_PIPETX5DATA10 (PIPETX5DATA[10], PIPETX5DATA_OUT[10]);
  buf B_PIPETX5DATA11 (PIPETX5DATA[11], PIPETX5DATA_OUT[11]);
  buf B_PIPETX5DATA12 (PIPETX5DATA[12], PIPETX5DATA_OUT[12]);
  buf B_PIPETX5DATA13 (PIPETX5DATA[13], PIPETX5DATA_OUT[13]);
  buf B_PIPETX5DATA14 (PIPETX5DATA[14], PIPETX5DATA_OUT[14]);
  buf B_PIPETX5DATA15 (PIPETX5DATA[15], PIPETX5DATA_OUT[15]);
  buf B_PIPETX5DATA16 (PIPETX5DATA[16], PIPETX5DATA_OUT[16]);
  buf B_PIPETX5DATA17 (PIPETX5DATA[17], PIPETX5DATA_OUT[17]);
  buf B_PIPETX5DATA18 (PIPETX5DATA[18], PIPETX5DATA_OUT[18]);
  buf B_PIPETX5DATA19 (PIPETX5DATA[19], PIPETX5DATA_OUT[19]);
  buf B_PIPETX5DATA2 (PIPETX5DATA[2], PIPETX5DATA_OUT[2]);
  buf B_PIPETX5DATA20 (PIPETX5DATA[20], PIPETX5DATA_OUT[20]);
  buf B_PIPETX5DATA21 (PIPETX5DATA[21], PIPETX5DATA_OUT[21]);
  buf B_PIPETX5DATA22 (PIPETX5DATA[22], PIPETX5DATA_OUT[22]);
  buf B_PIPETX5DATA23 (PIPETX5DATA[23], PIPETX5DATA_OUT[23]);
  buf B_PIPETX5DATA24 (PIPETX5DATA[24], PIPETX5DATA_OUT[24]);
  buf B_PIPETX5DATA25 (PIPETX5DATA[25], PIPETX5DATA_OUT[25]);
  buf B_PIPETX5DATA26 (PIPETX5DATA[26], PIPETX5DATA_OUT[26]);
  buf B_PIPETX5DATA27 (PIPETX5DATA[27], PIPETX5DATA_OUT[27]);
  buf B_PIPETX5DATA28 (PIPETX5DATA[28], PIPETX5DATA_OUT[28]);
  buf B_PIPETX5DATA29 (PIPETX5DATA[29], PIPETX5DATA_OUT[29]);
  buf B_PIPETX5DATA3 (PIPETX5DATA[3], PIPETX5DATA_OUT[3]);
  buf B_PIPETX5DATA30 (PIPETX5DATA[30], PIPETX5DATA_OUT[30]);
  buf B_PIPETX5DATA31 (PIPETX5DATA[31], PIPETX5DATA_OUT[31]);
  buf B_PIPETX5DATA4 (PIPETX5DATA[4], PIPETX5DATA_OUT[4]);
  buf B_PIPETX5DATA5 (PIPETX5DATA[5], PIPETX5DATA_OUT[5]);
  buf B_PIPETX5DATA6 (PIPETX5DATA[6], PIPETX5DATA_OUT[6]);
  buf B_PIPETX5DATA7 (PIPETX5DATA[7], PIPETX5DATA_OUT[7]);
  buf B_PIPETX5DATA8 (PIPETX5DATA[8], PIPETX5DATA_OUT[8]);
  buf B_PIPETX5DATA9 (PIPETX5DATA[9], PIPETX5DATA_OUT[9]);
  buf B_PIPETX5DATAVALID (PIPETX5DATAVALID, PIPETX5DATAVALID_OUT);
  buf B_PIPETX5ELECIDLE (PIPETX5ELECIDLE, PIPETX5ELECIDLE_OUT);
  buf B_PIPETX5EQCONTROL0 (PIPETX5EQCONTROL[0], PIPETX5EQCONTROL_OUT[0]);
  buf B_PIPETX5EQCONTROL1 (PIPETX5EQCONTROL[1], PIPETX5EQCONTROL_OUT[1]);
  buf B_PIPETX5EQDEEMPH0 (PIPETX5EQDEEMPH[0], PIPETX5EQDEEMPH_OUT[0]);
  buf B_PIPETX5EQDEEMPH1 (PIPETX5EQDEEMPH[1], PIPETX5EQDEEMPH_OUT[1]);
  buf B_PIPETX5EQDEEMPH2 (PIPETX5EQDEEMPH[2], PIPETX5EQDEEMPH_OUT[2]);
  buf B_PIPETX5EQDEEMPH3 (PIPETX5EQDEEMPH[3], PIPETX5EQDEEMPH_OUT[3]);
  buf B_PIPETX5EQDEEMPH4 (PIPETX5EQDEEMPH[4], PIPETX5EQDEEMPH_OUT[4]);
  buf B_PIPETX5EQDEEMPH5 (PIPETX5EQDEEMPH[5], PIPETX5EQDEEMPH_OUT[5]);
  buf B_PIPETX5EQPRESET0 (PIPETX5EQPRESET[0], PIPETX5EQPRESET_OUT[0]);
  buf B_PIPETX5EQPRESET1 (PIPETX5EQPRESET[1], PIPETX5EQPRESET_OUT[1]);
  buf B_PIPETX5EQPRESET2 (PIPETX5EQPRESET[2], PIPETX5EQPRESET_OUT[2]);
  buf B_PIPETX5EQPRESET3 (PIPETX5EQPRESET[3], PIPETX5EQPRESET_OUT[3]);
  buf B_PIPETX5POWERDOWN0 (PIPETX5POWERDOWN[0], PIPETX5POWERDOWN_OUT[0]);
  buf B_PIPETX5POWERDOWN1 (PIPETX5POWERDOWN[1], PIPETX5POWERDOWN_OUT[1]);
  buf B_PIPETX5STARTBLOCK (PIPETX5STARTBLOCK, PIPETX5STARTBLOCK_OUT);
  buf B_PIPETX5SYNCHEADER0 (PIPETX5SYNCHEADER[0], PIPETX5SYNCHEADER_OUT[0]);
  buf B_PIPETX5SYNCHEADER1 (PIPETX5SYNCHEADER[1], PIPETX5SYNCHEADER_OUT[1]);
  buf B_PIPETX6CHARISK0 (PIPETX6CHARISK[0], PIPETX6CHARISK_OUT[0]);
  buf B_PIPETX6CHARISK1 (PIPETX6CHARISK[1], PIPETX6CHARISK_OUT[1]);
  buf B_PIPETX6COMPLIANCE (PIPETX6COMPLIANCE, PIPETX6COMPLIANCE_OUT);
  buf B_PIPETX6DATA0 (PIPETX6DATA[0], PIPETX6DATA_OUT[0]);
  buf B_PIPETX6DATA1 (PIPETX6DATA[1], PIPETX6DATA_OUT[1]);
  buf B_PIPETX6DATA10 (PIPETX6DATA[10], PIPETX6DATA_OUT[10]);
  buf B_PIPETX6DATA11 (PIPETX6DATA[11], PIPETX6DATA_OUT[11]);
  buf B_PIPETX6DATA12 (PIPETX6DATA[12], PIPETX6DATA_OUT[12]);
  buf B_PIPETX6DATA13 (PIPETX6DATA[13], PIPETX6DATA_OUT[13]);
  buf B_PIPETX6DATA14 (PIPETX6DATA[14], PIPETX6DATA_OUT[14]);
  buf B_PIPETX6DATA15 (PIPETX6DATA[15], PIPETX6DATA_OUT[15]);
  buf B_PIPETX6DATA16 (PIPETX6DATA[16], PIPETX6DATA_OUT[16]);
  buf B_PIPETX6DATA17 (PIPETX6DATA[17], PIPETX6DATA_OUT[17]);
  buf B_PIPETX6DATA18 (PIPETX6DATA[18], PIPETX6DATA_OUT[18]);
  buf B_PIPETX6DATA19 (PIPETX6DATA[19], PIPETX6DATA_OUT[19]);
  buf B_PIPETX6DATA2 (PIPETX6DATA[2], PIPETX6DATA_OUT[2]);
  buf B_PIPETX6DATA20 (PIPETX6DATA[20], PIPETX6DATA_OUT[20]);
  buf B_PIPETX6DATA21 (PIPETX6DATA[21], PIPETX6DATA_OUT[21]);
  buf B_PIPETX6DATA22 (PIPETX6DATA[22], PIPETX6DATA_OUT[22]);
  buf B_PIPETX6DATA23 (PIPETX6DATA[23], PIPETX6DATA_OUT[23]);
  buf B_PIPETX6DATA24 (PIPETX6DATA[24], PIPETX6DATA_OUT[24]);
  buf B_PIPETX6DATA25 (PIPETX6DATA[25], PIPETX6DATA_OUT[25]);
  buf B_PIPETX6DATA26 (PIPETX6DATA[26], PIPETX6DATA_OUT[26]);
  buf B_PIPETX6DATA27 (PIPETX6DATA[27], PIPETX6DATA_OUT[27]);
  buf B_PIPETX6DATA28 (PIPETX6DATA[28], PIPETX6DATA_OUT[28]);
  buf B_PIPETX6DATA29 (PIPETX6DATA[29], PIPETX6DATA_OUT[29]);
  buf B_PIPETX6DATA3 (PIPETX6DATA[3], PIPETX6DATA_OUT[3]);
  buf B_PIPETX6DATA30 (PIPETX6DATA[30], PIPETX6DATA_OUT[30]);
  buf B_PIPETX6DATA31 (PIPETX6DATA[31], PIPETX6DATA_OUT[31]);
  buf B_PIPETX6DATA4 (PIPETX6DATA[4], PIPETX6DATA_OUT[4]);
  buf B_PIPETX6DATA5 (PIPETX6DATA[5], PIPETX6DATA_OUT[5]);
  buf B_PIPETX6DATA6 (PIPETX6DATA[6], PIPETX6DATA_OUT[6]);
  buf B_PIPETX6DATA7 (PIPETX6DATA[7], PIPETX6DATA_OUT[7]);
  buf B_PIPETX6DATA8 (PIPETX6DATA[8], PIPETX6DATA_OUT[8]);
  buf B_PIPETX6DATA9 (PIPETX6DATA[9], PIPETX6DATA_OUT[9]);
  buf B_PIPETX6DATAVALID (PIPETX6DATAVALID, PIPETX6DATAVALID_OUT);
  buf B_PIPETX6ELECIDLE (PIPETX6ELECIDLE, PIPETX6ELECIDLE_OUT);
  buf B_PIPETX6EQCONTROL0 (PIPETX6EQCONTROL[0], PIPETX6EQCONTROL_OUT[0]);
  buf B_PIPETX6EQCONTROL1 (PIPETX6EQCONTROL[1], PIPETX6EQCONTROL_OUT[1]);
  buf B_PIPETX6EQDEEMPH0 (PIPETX6EQDEEMPH[0], PIPETX6EQDEEMPH_OUT[0]);
  buf B_PIPETX6EQDEEMPH1 (PIPETX6EQDEEMPH[1], PIPETX6EQDEEMPH_OUT[1]);
  buf B_PIPETX6EQDEEMPH2 (PIPETX6EQDEEMPH[2], PIPETX6EQDEEMPH_OUT[2]);
  buf B_PIPETX6EQDEEMPH3 (PIPETX6EQDEEMPH[3], PIPETX6EQDEEMPH_OUT[3]);
  buf B_PIPETX6EQDEEMPH4 (PIPETX6EQDEEMPH[4], PIPETX6EQDEEMPH_OUT[4]);
  buf B_PIPETX6EQDEEMPH5 (PIPETX6EQDEEMPH[5], PIPETX6EQDEEMPH_OUT[5]);
  buf B_PIPETX6EQPRESET0 (PIPETX6EQPRESET[0], PIPETX6EQPRESET_OUT[0]);
  buf B_PIPETX6EQPRESET1 (PIPETX6EQPRESET[1], PIPETX6EQPRESET_OUT[1]);
  buf B_PIPETX6EQPRESET2 (PIPETX6EQPRESET[2], PIPETX6EQPRESET_OUT[2]);
  buf B_PIPETX6EQPRESET3 (PIPETX6EQPRESET[3], PIPETX6EQPRESET_OUT[3]);
  buf B_PIPETX6POWERDOWN0 (PIPETX6POWERDOWN[0], PIPETX6POWERDOWN_OUT[0]);
  buf B_PIPETX6POWERDOWN1 (PIPETX6POWERDOWN[1], PIPETX6POWERDOWN_OUT[1]);
  buf B_PIPETX6STARTBLOCK (PIPETX6STARTBLOCK, PIPETX6STARTBLOCK_OUT);
  buf B_PIPETX6SYNCHEADER0 (PIPETX6SYNCHEADER[0], PIPETX6SYNCHEADER_OUT[0]);
  buf B_PIPETX6SYNCHEADER1 (PIPETX6SYNCHEADER[1], PIPETX6SYNCHEADER_OUT[1]);
  buf B_PIPETX7CHARISK0 (PIPETX7CHARISK[0], PIPETX7CHARISK_OUT[0]);
  buf B_PIPETX7CHARISK1 (PIPETX7CHARISK[1], PIPETX7CHARISK_OUT[1]);
  buf B_PIPETX7COMPLIANCE (PIPETX7COMPLIANCE, PIPETX7COMPLIANCE_OUT);
  buf B_PIPETX7DATA0 (PIPETX7DATA[0], PIPETX7DATA_OUT[0]);
  buf B_PIPETX7DATA1 (PIPETX7DATA[1], PIPETX7DATA_OUT[1]);
  buf B_PIPETX7DATA10 (PIPETX7DATA[10], PIPETX7DATA_OUT[10]);
  buf B_PIPETX7DATA11 (PIPETX7DATA[11], PIPETX7DATA_OUT[11]);
  buf B_PIPETX7DATA12 (PIPETX7DATA[12], PIPETX7DATA_OUT[12]);
  buf B_PIPETX7DATA13 (PIPETX7DATA[13], PIPETX7DATA_OUT[13]);
  buf B_PIPETX7DATA14 (PIPETX7DATA[14], PIPETX7DATA_OUT[14]);
  buf B_PIPETX7DATA15 (PIPETX7DATA[15], PIPETX7DATA_OUT[15]);
  buf B_PIPETX7DATA16 (PIPETX7DATA[16], PIPETX7DATA_OUT[16]);
  buf B_PIPETX7DATA17 (PIPETX7DATA[17], PIPETX7DATA_OUT[17]);
  buf B_PIPETX7DATA18 (PIPETX7DATA[18], PIPETX7DATA_OUT[18]);
  buf B_PIPETX7DATA19 (PIPETX7DATA[19], PIPETX7DATA_OUT[19]);
  buf B_PIPETX7DATA2 (PIPETX7DATA[2], PIPETX7DATA_OUT[2]);
  buf B_PIPETX7DATA20 (PIPETX7DATA[20], PIPETX7DATA_OUT[20]);
  buf B_PIPETX7DATA21 (PIPETX7DATA[21], PIPETX7DATA_OUT[21]);
  buf B_PIPETX7DATA22 (PIPETX7DATA[22], PIPETX7DATA_OUT[22]);
  buf B_PIPETX7DATA23 (PIPETX7DATA[23], PIPETX7DATA_OUT[23]);
  buf B_PIPETX7DATA24 (PIPETX7DATA[24], PIPETX7DATA_OUT[24]);
  buf B_PIPETX7DATA25 (PIPETX7DATA[25], PIPETX7DATA_OUT[25]);
  buf B_PIPETX7DATA26 (PIPETX7DATA[26], PIPETX7DATA_OUT[26]);
  buf B_PIPETX7DATA27 (PIPETX7DATA[27], PIPETX7DATA_OUT[27]);
  buf B_PIPETX7DATA28 (PIPETX7DATA[28], PIPETX7DATA_OUT[28]);
  buf B_PIPETX7DATA29 (PIPETX7DATA[29], PIPETX7DATA_OUT[29]);
  buf B_PIPETX7DATA3 (PIPETX7DATA[3], PIPETX7DATA_OUT[3]);
  buf B_PIPETX7DATA30 (PIPETX7DATA[30], PIPETX7DATA_OUT[30]);
  buf B_PIPETX7DATA31 (PIPETX7DATA[31], PIPETX7DATA_OUT[31]);
  buf B_PIPETX7DATA4 (PIPETX7DATA[4], PIPETX7DATA_OUT[4]);
  buf B_PIPETX7DATA5 (PIPETX7DATA[5], PIPETX7DATA_OUT[5]);
  buf B_PIPETX7DATA6 (PIPETX7DATA[6], PIPETX7DATA_OUT[6]);
  buf B_PIPETX7DATA7 (PIPETX7DATA[7], PIPETX7DATA_OUT[7]);
  buf B_PIPETX7DATA8 (PIPETX7DATA[8], PIPETX7DATA_OUT[8]);
  buf B_PIPETX7DATA9 (PIPETX7DATA[9], PIPETX7DATA_OUT[9]);
  buf B_PIPETX7DATAVALID (PIPETX7DATAVALID, PIPETX7DATAVALID_OUT);
  buf B_PIPETX7ELECIDLE (PIPETX7ELECIDLE, PIPETX7ELECIDLE_OUT);
  buf B_PIPETX7EQCONTROL0 (PIPETX7EQCONTROL[0], PIPETX7EQCONTROL_OUT[0]);
  buf B_PIPETX7EQCONTROL1 (PIPETX7EQCONTROL[1], PIPETX7EQCONTROL_OUT[1]);
  buf B_PIPETX7EQDEEMPH0 (PIPETX7EQDEEMPH[0], PIPETX7EQDEEMPH_OUT[0]);
  buf B_PIPETX7EQDEEMPH1 (PIPETX7EQDEEMPH[1], PIPETX7EQDEEMPH_OUT[1]);
  buf B_PIPETX7EQDEEMPH2 (PIPETX7EQDEEMPH[2], PIPETX7EQDEEMPH_OUT[2]);
  buf B_PIPETX7EQDEEMPH3 (PIPETX7EQDEEMPH[3], PIPETX7EQDEEMPH_OUT[3]);
  buf B_PIPETX7EQDEEMPH4 (PIPETX7EQDEEMPH[4], PIPETX7EQDEEMPH_OUT[4]);
  buf B_PIPETX7EQDEEMPH5 (PIPETX7EQDEEMPH[5], PIPETX7EQDEEMPH_OUT[5]);
  buf B_PIPETX7EQPRESET0 (PIPETX7EQPRESET[0], PIPETX7EQPRESET_OUT[0]);
  buf B_PIPETX7EQPRESET1 (PIPETX7EQPRESET[1], PIPETX7EQPRESET_OUT[1]);
  buf B_PIPETX7EQPRESET2 (PIPETX7EQPRESET[2], PIPETX7EQPRESET_OUT[2]);
  buf B_PIPETX7EQPRESET3 (PIPETX7EQPRESET[3], PIPETX7EQPRESET_OUT[3]);
  buf B_PIPETX7POWERDOWN0 (PIPETX7POWERDOWN[0], PIPETX7POWERDOWN_OUT[0]);
  buf B_PIPETX7POWERDOWN1 (PIPETX7POWERDOWN[1], PIPETX7POWERDOWN_OUT[1]);
  buf B_PIPETX7STARTBLOCK (PIPETX7STARTBLOCK, PIPETX7STARTBLOCK_OUT);
  buf B_PIPETX7SYNCHEADER0 (PIPETX7SYNCHEADER[0], PIPETX7SYNCHEADER_OUT[0]);
  buf B_PIPETX7SYNCHEADER1 (PIPETX7SYNCHEADER[1], PIPETX7SYNCHEADER_OUT[1]);
  buf B_PIPETXDEEMPH (PIPETXDEEMPH, PIPETXDEEMPH_OUT);
  buf B_PIPETXMARGIN0 (PIPETXMARGIN[0], PIPETXMARGIN_OUT[0]);
  buf B_PIPETXMARGIN1 (PIPETXMARGIN[1], PIPETXMARGIN_OUT[1]);
  buf B_PIPETXMARGIN2 (PIPETXMARGIN[2], PIPETXMARGIN_OUT[2]);
  buf B_PIPETXRATE0 (PIPETXRATE[0], PIPETXRATE_OUT[0]);
  buf B_PIPETXRATE1 (PIPETXRATE[1], PIPETXRATE_OUT[1]);
  buf B_PIPETXRCVRDET (PIPETXRCVRDET, PIPETXRCVRDET_OUT);
  buf B_PIPETXRESET (PIPETXRESET, PIPETXRESET_OUT);
  buf B_PIPETXSWING (PIPETXSWING, PIPETXSWING_OUT);
  buf B_PLEQINPROGRESS (PLEQINPROGRESS, PLEQINPROGRESS_OUT);
  buf B_PLEQPHASE0 (PLEQPHASE[0], PLEQPHASE_OUT[0]);
  buf B_PLEQPHASE1 (PLEQPHASE[1], PLEQPHASE_OUT[1]);
  buf B_PLGEN3PCSRXSLIDE0 (PLGEN3PCSRXSLIDE[0], PLGEN3PCSRXSLIDE_OUT[0]);
  buf B_PLGEN3PCSRXSLIDE1 (PLGEN3PCSRXSLIDE[1], PLGEN3PCSRXSLIDE_OUT[1]);
  buf B_PLGEN3PCSRXSLIDE2 (PLGEN3PCSRXSLIDE[2], PLGEN3PCSRXSLIDE_OUT[2]);
  buf B_PLGEN3PCSRXSLIDE3 (PLGEN3PCSRXSLIDE[3], PLGEN3PCSRXSLIDE_OUT[3]);
  buf B_PLGEN3PCSRXSLIDE4 (PLGEN3PCSRXSLIDE[4], PLGEN3PCSRXSLIDE_OUT[4]);
  buf B_PLGEN3PCSRXSLIDE5 (PLGEN3PCSRXSLIDE[5], PLGEN3PCSRXSLIDE_OUT[5]);
  buf B_PLGEN3PCSRXSLIDE6 (PLGEN3PCSRXSLIDE[6], PLGEN3PCSRXSLIDE_OUT[6]);
  buf B_PLGEN3PCSRXSLIDE7 (PLGEN3PCSRXSLIDE[7], PLGEN3PCSRXSLIDE_OUT[7]);
  buf B_SAXISCCTREADY0 (SAXISCCTREADY[0], SAXISCCTREADY_OUT[0]);
  buf B_SAXISCCTREADY1 (SAXISCCTREADY[1], SAXISCCTREADY_OUT[1]);
  buf B_SAXISCCTREADY2 (SAXISCCTREADY[2], SAXISCCTREADY_OUT[2]);
  buf B_SAXISCCTREADY3 (SAXISCCTREADY[3], SAXISCCTREADY_OUT[3]);
  buf B_SAXISRQTREADY0 (SAXISRQTREADY[0], SAXISRQTREADY_OUT[0]);
  buf B_SAXISRQTREADY1 (SAXISRQTREADY[1], SAXISRQTREADY_OUT[1]);
  buf B_SAXISRQTREADY2 (SAXISRQTREADY[2], SAXISRQTREADY_OUT[2]);
  buf B_SAXISRQTREADY3 (SAXISRQTREADY[3], SAXISRQTREADY_OUT[3]);

  buf B_CFGCONFIGSPACEENABLE (CFGCONFIGSPACEENABLE_IN, CFGCONFIGSPACEENABLE);
  buf B_CFGDEVID0 (CFGDEVID_IN[0], CFGDEVID[0]);
  buf B_CFGDEVID1 (CFGDEVID_IN[1], CFGDEVID[1]);
  buf B_CFGDEVID10 (CFGDEVID_IN[10], CFGDEVID[10]);
  buf B_CFGDEVID11 (CFGDEVID_IN[11], CFGDEVID[11]);
  buf B_CFGDEVID12 (CFGDEVID_IN[12], CFGDEVID[12]);
  buf B_CFGDEVID13 (CFGDEVID_IN[13], CFGDEVID[13]);
  buf B_CFGDEVID14 (CFGDEVID_IN[14], CFGDEVID[14]);
  buf B_CFGDEVID15 (CFGDEVID_IN[15], CFGDEVID[15]);
  buf B_CFGDEVID2 (CFGDEVID_IN[2], CFGDEVID[2]);
  buf B_CFGDEVID3 (CFGDEVID_IN[3], CFGDEVID[3]);
  buf B_CFGDEVID4 (CFGDEVID_IN[4], CFGDEVID[4]);
  buf B_CFGDEVID5 (CFGDEVID_IN[5], CFGDEVID[5]);
  buf B_CFGDEVID6 (CFGDEVID_IN[6], CFGDEVID[6]);
  buf B_CFGDEVID7 (CFGDEVID_IN[7], CFGDEVID[7]);
  buf B_CFGDEVID8 (CFGDEVID_IN[8], CFGDEVID[8]);
  buf B_CFGDEVID9 (CFGDEVID_IN[9], CFGDEVID[9]);
  buf B_CFGDSBUSNUMBER0 (CFGDSBUSNUMBER_IN[0], CFGDSBUSNUMBER[0]);
  buf B_CFGDSBUSNUMBER1 (CFGDSBUSNUMBER_IN[1], CFGDSBUSNUMBER[1]);
  buf B_CFGDSBUSNUMBER2 (CFGDSBUSNUMBER_IN[2], CFGDSBUSNUMBER[2]);
  buf B_CFGDSBUSNUMBER3 (CFGDSBUSNUMBER_IN[3], CFGDSBUSNUMBER[3]);
  buf B_CFGDSBUSNUMBER4 (CFGDSBUSNUMBER_IN[4], CFGDSBUSNUMBER[4]);
  buf B_CFGDSBUSNUMBER5 (CFGDSBUSNUMBER_IN[5], CFGDSBUSNUMBER[5]);
  buf B_CFGDSBUSNUMBER6 (CFGDSBUSNUMBER_IN[6], CFGDSBUSNUMBER[6]);
  buf B_CFGDSBUSNUMBER7 (CFGDSBUSNUMBER_IN[7], CFGDSBUSNUMBER[7]);
  buf B_CFGDSDEVICENUMBER0 (CFGDSDEVICENUMBER_IN[0], CFGDSDEVICENUMBER[0]);
  buf B_CFGDSDEVICENUMBER1 (CFGDSDEVICENUMBER_IN[1], CFGDSDEVICENUMBER[1]);
  buf B_CFGDSDEVICENUMBER2 (CFGDSDEVICENUMBER_IN[2], CFGDSDEVICENUMBER[2]);
  buf B_CFGDSDEVICENUMBER3 (CFGDSDEVICENUMBER_IN[3], CFGDSDEVICENUMBER[3]);
  buf B_CFGDSDEVICENUMBER4 (CFGDSDEVICENUMBER_IN[4], CFGDSDEVICENUMBER[4]);
  buf B_CFGDSFUNCTIONNUMBER0 (CFGDSFUNCTIONNUMBER_IN[0], CFGDSFUNCTIONNUMBER[0]);
  buf B_CFGDSFUNCTIONNUMBER1 (CFGDSFUNCTIONNUMBER_IN[1], CFGDSFUNCTIONNUMBER[1]);
  buf B_CFGDSFUNCTIONNUMBER2 (CFGDSFUNCTIONNUMBER_IN[2], CFGDSFUNCTIONNUMBER[2]);
  buf B_CFGDSN0 (CFGDSN_IN[0], CFGDSN[0]);
  buf B_CFGDSN1 (CFGDSN_IN[1], CFGDSN[1]);
  buf B_CFGDSN10 (CFGDSN_IN[10], CFGDSN[10]);
  buf B_CFGDSN11 (CFGDSN_IN[11], CFGDSN[11]);
  buf B_CFGDSN12 (CFGDSN_IN[12], CFGDSN[12]);
  buf B_CFGDSN13 (CFGDSN_IN[13], CFGDSN[13]);
  buf B_CFGDSN14 (CFGDSN_IN[14], CFGDSN[14]);
  buf B_CFGDSN15 (CFGDSN_IN[15], CFGDSN[15]);
  buf B_CFGDSN16 (CFGDSN_IN[16], CFGDSN[16]);
  buf B_CFGDSN17 (CFGDSN_IN[17], CFGDSN[17]);
  buf B_CFGDSN18 (CFGDSN_IN[18], CFGDSN[18]);
  buf B_CFGDSN19 (CFGDSN_IN[19], CFGDSN[19]);
  buf B_CFGDSN2 (CFGDSN_IN[2], CFGDSN[2]);
  buf B_CFGDSN20 (CFGDSN_IN[20], CFGDSN[20]);
  buf B_CFGDSN21 (CFGDSN_IN[21], CFGDSN[21]);
  buf B_CFGDSN22 (CFGDSN_IN[22], CFGDSN[22]);
  buf B_CFGDSN23 (CFGDSN_IN[23], CFGDSN[23]);
  buf B_CFGDSN24 (CFGDSN_IN[24], CFGDSN[24]);
  buf B_CFGDSN25 (CFGDSN_IN[25], CFGDSN[25]);
  buf B_CFGDSN26 (CFGDSN_IN[26], CFGDSN[26]);
  buf B_CFGDSN27 (CFGDSN_IN[27], CFGDSN[27]);
  buf B_CFGDSN28 (CFGDSN_IN[28], CFGDSN[28]);
  buf B_CFGDSN29 (CFGDSN_IN[29], CFGDSN[29]);
  buf B_CFGDSN3 (CFGDSN_IN[3], CFGDSN[3]);
  buf B_CFGDSN30 (CFGDSN_IN[30], CFGDSN[30]);
  buf B_CFGDSN31 (CFGDSN_IN[31], CFGDSN[31]);
  buf B_CFGDSN32 (CFGDSN_IN[32], CFGDSN[32]);
  buf B_CFGDSN33 (CFGDSN_IN[33], CFGDSN[33]);
  buf B_CFGDSN34 (CFGDSN_IN[34], CFGDSN[34]);
  buf B_CFGDSN35 (CFGDSN_IN[35], CFGDSN[35]);
  buf B_CFGDSN36 (CFGDSN_IN[36], CFGDSN[36]);
  buf B_CFGDSN37 (CFGDSN_IN[37], CFGDSN[37]);
  buf B_CFGDSN38 (CFGDSN_IN[38], CFGDSN[38]);
  buf B_CFGDSN39 (CFGDSN_IN[39], CFGDSN[39]);
  buf B_CFGDSN4 (CFGDSN_IN[4], CFGDSN[4]);
  buf B_CFGDSN40 (CFGDSN_IN[40], CFGDSN[40]);
  buf B_CFGDSN41 (CFGDSN_IN[41], CFGDSN[41]);
  buf B_CFGDSN42 (CFGDSN_IN[42], CFGDSN[42]);
  buf B_CFGDSN43 (CFGDSN_IN[43], CFGDSN[43]);
  buf B_CFGDSN44 (CFGDSN_IN[44], CFGDSN[44]);
  buf B_CFGDSN45 (CFGDSN_IN[45], CFGDSN[45]);
  buf B_CFGDSN46 (CFGDSN_IN[46], CFGDSN[46]);
  buf B_CFGDSN47 (CFGDSN_IN[47], CFGDSN[47]);
  buf B_CFGDSN48 (CFGDSN_IN[48], CFGDSN[48]);
  buf B_CFGDSN49 (CFGDSN_IN[49], CFGDSN[49]);
  buf B_CFGDSN5 (CFGDSN_IN[5], CFGDSN[5]);
  buf B_CFGDSN50 (CFGDSN_IN[50], CFGDSN[50]);
  buf B_CFGDSN51 (CFGDSN_IN[51], CFGDSN[51]);
  buf B_CFGDSN52 (CFGDSN_IN[52], CFGDSN[52]);
  buf B_CFGDSN53 (CFGDSN_IN[53], CFGDSN[53]);
  buf B_CFGDSN54 (CFGDSN_IN[54], CFGDSN[54]);
  buf B_CFGDSN55 (CFGDSN_IN[55], CFGDSN[55]);
  buf B_CFGDSN56 (CFGDSN_IN[56], CFGDSN[56]);
  buf B_CFGDSN57 (CFGDSN_IN[57], CFGDSN[57]);
  buf B_CFGDSN58 (CFGDSN_IN[58], CFGDSN[58]);
  buf B_CFGDSN59 (CFGDSN_IN[59], CFGDSN[59]);
  buf B_CFGDSN6 (CFGDSN_IN[6], CFGDSN[6]);
  buf B_CFGDSN60 (CFGDSN_IN[60], CFGDSN[60]);
  buf B_CFGDSN61 (CFGDSN_IN[61], CFGDSN[61]);
  buf B_CFGDSN62 (CFGDSN_IN[62], CFGDSN[62]);
  buf B_CFGDSN63 (CFGDSN_IN[63], CFGDSN[63]);
  buf B_CFGDSN7 (CFGDSN_IN[7], CFGDSN[7]);
  buf B_CFGDSN8 (CFGDSN_IN[8], CFGDSN[8]);
  buf B_CFGDSN9 (CFGDSN_IN[9], CFGDSN[9]);
  buf B_CFGDSPORTNUMBER0 (CFGDSPORTNUMBER_IN[0], CFGDSPORTNUMBER[0]);
  buf B_CFGDSPORTNUMBER1 (CFGDSPORTNUMBER_IN[1], CFGDSPORTNUMBER[1]);
  buf B_CFGDSPORTNUMBER2 (CFGDSPORTNUMBER_IN[2], CFGDSPORTNUMBER[2]);
  buf B_CFGDSPORTNUMBER3 (CFGDSPORTNUMBER_IN[3], CFGDSPORTNUMBER[3]);
  buf B_CFGDSPORTNUMBER4 (CFGDSPORTNUMBER_IN[4], CFGDSPORTNUMBER[4]);
  buf B_CFGDSPORTNUMBER5 (CFGDSPORTNUMBER_IN[5], CFGDSPORTNUMBER[5]);
  buf B_CFGDSPORTNUMBER6 (CFGDSPORTNUMBER_IN[6], CFGDSPORTNUMBER[6]);
  buf B_CFGDSPORTNUMBER7 (CFGDSPORTNUMBER_IN[7], CFGDSPORTNUMBER[7]);
  buf B_CFGERRCORIN (CFGERRCORIN_IN, CFGERRCORIN);
  buf B_CFGERRUNCORIN (CFGERRUNCORIN_IN, CFGERRUNCORIN);
  buf B_CFGEXTREADDATA0 (CFGEXTREADDATA_IN[0], CFGEXTREADDATA[0]);
  buf B_CFGEXTREADDATA1 (CFGEXTREADDATA_IN[1], CFGEXTREADDATA[1]);
  buf B_CFGEXTREADDATA10 (CFGEXTREADDATA_IN[10], CFGEXTREADDATA[10]);
  buf B_CFGEXTREADDATA11 (CFGEXTREADDATA_IN[11], CFGEXTREADDATA[11]);
  buf B_CFGEXTREADDATA12 (CFGEXTREADDATA_IN[12], CFGEXTREADDATA[12]);
  buf B_CFGEXTREADDATA13 (CFGEXTREADDATA_IN[13], CFGEXTREADDATA[13]);
  buf B_CFGEXTREADDATA14 (CFGEXTREADDATA_IN[14], CFGEXTREADDATA[14]);
  buf B_CFGEXTREADDATA15 (CFGEXTREADDATA_IN[15], CFGEXTREADDATA[15]);
  buf B_CFGEXTREADDATA16 (CFGEXTREADDATA_IN[16], CFGEXTREADDATA[16]);
  buf B_CFGEXTREADDATA17 (CFGEXTREADDATA_IN[17], CFGEXTREADDATA[17]);
  buf B_CFGEXTREADDATA18 (CFGEXTREADDATA_IN[18], CFGEXTREADDATA[18]);
  buf B_CFGEXTREADDATA19 (CFGEXTREADDATA_IN[19], CFGEXTREADDATA[19]);
  buf B_CFGEXTREADDATA2 (CFGEXTREADDATA_IN[2], CFGEXTREADDATA[2]);
  buf B_CFGEXTREADDATA20 (CFGEXTREADDATA_IN[20], CFGEXTREADDATA[20]);
  buf B_CFGEXTREADDATA21 (CFGEXTREADDATA_IN[21], CFGEXTREADDATA[21]);
  buf B_CFGEXTREADDATA22 (CFGEXTREADDATA_IN[22], CFGEXTREADDATA[22]);
  buf B_CFGEXTREADDATA23 (CFGEXTREADDATA_IN[23], CFGEXTREADDATA[23]);
  buf B_CFGEXTREADDATA24 (CFGEXTREADDATA_IN[24], CFGEXTREADDATA[24]);
  buf B_CFGEXTREADDATA25 (CFGEXTREADDATA_IN[25], CFGEXTREADDATA[25]);
  buf B_CFGEXTREADDATA26 (CFGEXTREADDATA_IN[26], CFGEXTREADDATA[26]);
  buf B_CFGEXTREADDATA27 (CFGEXTREADDATA_IN[27], CFGEXTREADDATA[27]);
  buf B_CFGEXTREADDATA28 (CFGEXTREADDATA_IN[28], CFGEXTREADDATA[28]);
  buf B_CFGEXTREADDATA29 (CFGEXTREADDATA_IN[29], CFGEXTREADDATA[29]);
  buf B_CFGEXTREADDATA3 (CFGEXTREADDATA_IN[3], CFGEXTREADDATA[3]);
  buf B_CFGEXTREADDATA30 (CFGEXTREADDATA_IN[30], CFGEXTREADDATA[30]);
  buf B_CFGEXTREADDATA31 (CFGEXTREADDATA_IN[31], CFGEXTREADDATA[31]);
  buf B_CFGEXTREADDATA4 (CFGEXTREADDATA_IN[4], CFGEXTREADDATA[4]);
  buf B_CFGEXTREADDATA5 (CFGEXTREADDATA_IN[5], CFGEXTREADDATA[5]);
  buf B_CFGEXTREADDATA6 (CFGEXTREADDATA_IN[6], CFGEXTREADDATA[6]);
  buf B_CFGEXTREADDATA7 (CFGEXTREADDATA_IN[7], CFGEXTREADDATA[7]);
  buf B_CFGEXTREADDATA8 (CFGEXTREADDATA_IN[8], CFGEXTREADDATA[8]);
  buf B_CFGEXTREADDATA9 (CFGEXTREADDATA_IN[9], CFGEXTREADDATA[9]);
  buf B_CFGEXTREADDATAVALID (CFGEXTREADDATAVALID_IN, CFGEXTREADDATAVALID);
  buf B_CFGFCSEL0 (CFGFCSEL_IN[0], CFGFCSEL[0]);
  buf B_CFGFCSEL1 (CFGFCSEL_IN[1], CFGFCSEL[1]);
  buf B_CFGFCSEL2 (CFGFCSEL_IN[2], CFGFCSEL[2]);
  buf B_CFGFLRDONE0 (CFGFLRDONE_IN[0], CFGFLRDONE[0]);
  buf B_CFGFLRDONE1 (CFGFLRDONE_IN[1], CFGFLRDONE[1]);
  buf B_CFGHOTRESETIN (CFGHOTRESETIN_IN, CFGHOTRESETIN);
  buf B_CFGINPUTUPDATEREQUEST (CFGINPUTUPDATEREQUEST_IN, CFGINPUTUPDATEREQUEST);
  buf B_CFGINTERRUPTINT0 (CFGINTERRUPTINT_IN[0], CFGINTERRUPTINT[0]);
  buf B_CFGINTERRUPTINT1 (CFGINTERRUPTINT_IN[1], CFGINTERRUPTINT[1]);
  buf B_CFGINTERRUPTINT2 (CFGINTERRUPTINT_IN[2], CFGINTERRUPTINT[2]);
  buf B_CFGINTERRUPTINT3 (CFGINTERRUPTINT_IN[3], CFGINTERRUPTINT[3]);
  buf B_CFGINTERRUPTMSIATTR0 (CFGINTERRUPTMSIATTR_IN[0], CFGINTERRUPTMSIATTR[0]);
  buf B_CFGINTERRUPTMSIATTR1 (CFGINTERRUPTMSIATTR_IN[1], CFGINTERRUPTMSIATTR[1]);
  buf B_CFGINTERRUPTMSIATTR2 (CFGINTERRUPTMSIATTR_IN[2], CFGINTERRUPTMSIATTR[2]);
  buf B_CFGINTERRUPTMSIFUNCTIONNUMBER0 (CFGINTERRUPTMSIFUNCTIONNUMBER_IN[0], CFGINTERRUPTMSIFUNCTIONNUMBER[0]);
  buf B_CFGINTERRUPTMSIFUNCTIONNUMBER1 (CFGINTERRUPTMSIFUNCTIONNUMBER_IN[1], CFGINTERRUPTMSIFUNCTIONNUMBER[1]);
  buf B_CFGINTERRUPTMSIFUNCTIONNUMBER2 (CFGINTERRUPTMSIFUNCTIONNUMBER_IN[2], CFGINTERRUPTMSIFUNCTIONNUMBER[2]);
  buf B_CFGINTERRUPTMSIINT0 (CFGINTERRUPTMSIINT_IN[0], CFGINTERRUPTMSIINT[0]);
  buf B_CFGINTERRUPTMSIINT1 (CFGINTERRUPTMSIINT_IN[1], CFGINTERRUPTMSIINT[1]);
  buf B_CFGINTERRUPTMSIINT10 (CFGINTERRUPTMSIINT_IN[10], CFGINTERRUPTMSIINT[10]);
  buf B_CFGINTERRUPTMSIINT11 (CFGINTERRUPTMSIINT_IN[11], CFGINTERRUPTMSIINT[11]);
  buf B_CFGINTERRUPTMSIINT12 (CFGINTERRUPTMSIINT_IN[12], CFGINTERRUPTMSIINT[12]);
  buf B_CFGINTERRUPTMSIINT13 (CFGINTERRUPTMSIINT_IN[13], CFGINTERRUPTMSIINT[13]);
  buf B_CFGINTERRUPTMSIINT14 (CFGINTERRUPTMSIINT_IN[14], CFGINTERRUPTMSIINT[14]);
  buf B_CFGINTERRUPTMSIINT15 (CFGINTERRUPTMSIINT_IN[15], CFGINTERRUPTMSIINT[15]);
  buf B_CFGINTERRUPTMSIINT16 (CFGINTERRUPTMSIINT_IN[16], CFGINTERRUPTMSIINT[16]);
  buf B_CFGINTERRUPTMSIINT17 (CFGINTERRUPTMSIINT_IN[17], CFGINTERRUPTMSIINT[17]);
  buf B_CFGINTERRUPTMSIINT18 (CFGINTERRUPTMSIINT_IN[18], CFGINTERRUPTMSIINT[18]);
  buf B_CFGINTERRUPTMSIINT19 (CFGINTERRUPTMSIINT_IN[19], CFGINTERRUPTMSIINT[19]);
  buf B_CFGINTERRUPTMSIINT2 (CFGINTERRUPTMSIINT_IN[2], CFGINTERRUPTMSIINT[2]);
  buf B_CFGINTERRUPTMSIINT20 (CFGINTERRUPTMSIINT_IN[20], CFGINTERRUPTMSIINT[20]);
  buf B_CFGINTERRUPTMSIINT21 (CFGINTERRUPTMSIINT_IN[21], CFGINTERRUPTMSIINT[21]);
  buf B_CFGINTERRUPTMSIINT22 (CFGINTERRUPTMSIINT_IN[22], CFGINTERRUPTMSIINT[22]);
  buf B_CFGINTERRUPTMSIINT23 (CFGINTERRUPTMSIINT_IN[23], CFGINTERRUPTMSIINT[23]);
  buf B_CFGINTERRUPTMSIINT24 (CFGINTERRUPTMSIINT_IN[24], CFGINTERRUPTMSIINT[24]);
  buf B_CFGINTERRUPTMSIINT25 (CFGINTERRUPTMSIINT_IN[25], CFGINTERRUPTMSIINT[25]);
  buf B_CFGINTERRUPTMSIINT26 (CFGINTERRUPTMSIINT_IN[26], CFGINTERRUPTMSIINT[26]);
  buf B_CFGINTERRUPTMSIINT27 (CFGINTERRUPTMSIINT_IN[27], CFGINTERRUPTMSIINT[27]);
  buf B_CFGINTERRUPTMSIINT28 (CFGINTERRUPTMSIINT_IN[28], CFGINTERRUPTMSIINT[28]);
  buf B_CFGINTERRUPTMSIINT29 (CFGINTERRUPTMSIINT_IN[29], CFGINTERRUPTMSIINT[29]);
  buf B_CFGINTERRUPTMSIINT3 (CFGINTERRUPTMSIINT_IN[3], CFGINTERRUPTMSIINT[3]);
  buf B_CFGINTERRUPTMSIINT30 (CFGINTERRUPTMSIINT_IN[30], CFGINTERRUPTMSIINT[30]);
  buf B_CFGINTERRUPTMSIINT31 (CFGINTERRUPTMSIINT_IN[31], CFGINTERRUPTMSIINT[31]);
  buf B_CFGINTERRUPTMSIINT4 (CFGINTERRUPTMSIINT_IN[4], CFGINTERRUPTMSIINT[4]);
  buf B_CFGINTERRUPTMSIINT5 (CFGINTERRUPTMSIINT_IN[5], CFGINTERRUPTMSIINT[5]);
  buf B_CFGINTERRUPTMSIINT6 (CFGINTERRUPTMSIINT_IN[6], CFGINTERRUPTMSIINT[6]);
  buf B_CFGINTERRUPTMSIINT7 (CFGINTERRUPTMSIINT_IN[7], CFGINTERRUPTMSIINT[7]);
  buf B_CFGINTERRUPTMSIINT8 (CFGINTERRUPTMSIINT_IN[8], CFGINTERRUPTMSIINT[8]);
  buf B_CFGINTERRUPTMSIINT9 (CFGINTERRUPTMSIINT_IN[9], CFGINTERRUPTMSIINT[9]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS0 (CFGINTERRUPTMSIPENDINGSTATUS_IN[0], CFGINTERRUPTMSIPENDINGSTATUS[0]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS1 (CFGINTERRUPTMSIPENDINGSTATUS_IN[1], CFGINTERRUPTMSIPENDINGSTATUS[1]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS10 (CFGINTERRUPTMSIPENDINGSTATUS_IN[10], CFGINTERRUPTMSIPENDINGSTATUS[10]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS11 (CFGINTERRUPTMSIPENDINGSTATUS_IN[11], CFGINTERRUPTMSIPENDINGSTATUS[11]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS12 (CFGINTERRUPTMSIPENDINGSTATUS_IN[12], CFGINTERRUPTMSIPENDINGSTATUS[12]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS13 (CFGINTERRUPTMSIPENDINGSTATUS_IN[13], CFGINTERRUPTMSIPENDINGSTATUS[13]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS14 (CFGINTERRUPTMSIPENDINGSTATUS_IN[14], CFGINTERRUPTMSIPENDINGSTATUS[14]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS15 (CFGINTERRUPTMSIPENDINGSTATUS_IN[15], CFGINTERRUPTMSIPENDINGSTATUS[15]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS16 (CFGINTERRUPTMSIPENDINGSTATUS_IN[16], CFGINTERRUPTMSIPENDINGSTATUS[16]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS17 (CFGINTERRUPTMSIPENDINGSTATUS_IN[17], CFGINTERRUPTMSIPENDINGSTATUS[17]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS18 (CFGINTERRUPTMSIPENDINGSTATUS_IN[18], CFGINTERRUPTMSIPENDINGSTATUS[18]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS19 (CFGINTERRUPTMSIPENDINGSTATUS_IN[19], CFGINTERRUPTMSIPENDINGSTATUS[19]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS2 (CFGINTERRUPTMSIPENDINGSTATUS_IN[2], CFGINTERRUPTMSIPENDINGSTATUS[2]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS20 (CFGINTERRUPTMSIPENDINGSTATUS_IN[20], CFGINTERRUPTMSIPENDINGSTATUS[20]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS21 (CFGINTERRUPTMSIPENDINGSTATUS_IN[21], CFGINTERRUPTMSIPENDINGSTATUS[21]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS22 (CFGINTERRUPTMSIPENDINGSTATUS_IN[22], CFGINTERRUPTMSIPENDINGSTATUS[22]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS23 (CFGINTERRUPTMSIPENDINGSTATUS_IN[23], CFGINTERRUPTMSIPENDINGSTATUS[23]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS24 (CFGINTERRUPTMSIPENDINGSTATUS_IN[24], CFGINTERRUPTMSIPENDINGSTATUS[24]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS25 (CFGINTERRUPTMSIPENDINGSTATUS_IN[25], CFGINTERRUPTMSIPENDINGSTATUS[25]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS26 (CFGINTERRUPTMSIPENDINGSTATUS_IN[26], CFGINTERRUPTMSIPENDINGSTATUS[26]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS27 (CFGINTERRUPTMSIPENDINGSTATUS_IN[27], CFGINTERRUPTMSIPENDINGSTATUS[27]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS28 (CFGINTERRUPTMSIPENDINGSTATUS_IN[28], CFGINTERRUPTMSIPENDINGSTATUS[28]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS29 (CFGINTERRUPTMSIPENDINGSTATUS_IN[29], CFGINTERRUPTMSIPENDINGSTATUS[29]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS3 (CFGINTERRUPTMSIPENDINGSTATUS_IN[3], CFGINTERRUPTMSIPENDINGSTATUS[3]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS30 (CFGINTERRUPTMSIPENDINGSTATUS_IN[30], CFGINTERRUPTMSIPENDINGSTATUS[30]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS31 (CFGINTERRUPTMSIPENDINGSTATUS_IN[31], CFGINTERRUPTMSIPENDINGSTATUS[31]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS32 (CFGINTERRUPTMSIPENDINGSTATUS_IN[32], CFGINTERRUPTMSIPENDINGSTATUS[32]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS33 (CFGINTERRUPTMSIPENDINGSTATUS_IN[33], CFGINTERRUPTMSIPENDINGSTATUS[33]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS34 (CFGINTERRUPTMSIPENDINGSTATUS_IN[34], CFGINTERRUPTMSIPENDINGSTATUS[34]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS35 (CFGINTERRUPTMSIPENDINGSTATUS_IN[35], CFGINTERRUPTMSIPENDINGSTATUS[35]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS36 (CFGINTERRUPTMSIPENDINGSTATUS_IN[36], CFGINTERRUPTMSIPENDINGSTATUS[36]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS37 (CFGINTERRUPTMSIPENDINGSTATUS_IN[37], CFGINTERRUPTMSIPENDINGSTATUS[37]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS38 (CFGINTERRUPTMSIPENDINGSTATUS_IN[38], CFGINTERRUPTMSIPENDINGSTATUS[38]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS39 (CFGINTERRUPTMSIPENDINGSTATUS_IN[39], CFGINTERRUPTMSIPENDINGSTATUS[39]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS4 (CFGINTERRUPTMSIPENDINGSTATUS_IN[4], CFGINTERRUPTMSIPENDINGSTATUS[4]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS40 (CFGINTERRUPTMSIPENDINGSTATUS_IN[40], CFGINTERRUPTMSIPENDINGSTATUS[40]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS41 (CFGINTERRUPTMSIPENDINGSTATUS_IN[41], CFGINTERRUPTMSIPENDINGSTATUS[41]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS42 (CFGINTERRUPTMSIPENDINGSTATUS_IN[42], CFGINTERRUPTMSIPENDINGSTATUS[42]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS43 (CFGINTERRUPTMSIPENDINGSTATUS_IN[43], CFGINTERRUPTMSIPENDINGSTATUS[43]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS44 (CFGINTERRUPTMSIPENDINGSTATUS_IN[44], CFGINTERRUPTMSIPENDINGSTATUS[44]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS45 (CFGINTERRUPTMSIPENDINGSTATUS_IN[45], CFGINTERRUPTMSIPENDINGSTATUS[45]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS46 (CFGINTERRUPTMSIPENDINGSTATUS_IN[46], CFGINTERRUPTMSIPENDINGSTATUS[46]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS47 (CFGINTERRUPTMSIPENDINGSTATUS_IN[47], CFGINTERRUPTMSIPENDINGSTATUS[47]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS48 (CFGINTERRUPTMSIPENDINGSTATUS_IN[48], CFGINTERRUPTMSIPENDINGSTATUS[48]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS49 (CFGINTERRUPTMSIPENDINGSTATUS_IN[49], CFGINTERRUPTMSIPENDINGSTATUS[49]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS5 (CFGINTERRUPTMSIPENDINGSTATUS_IN[5], CFGINTERRUPTMSIPENDINGSTATUS[5]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS50 (CFGINTERRUPTMSIPENDINGSTATUS_IN[50], CFGINTERRUPTMSIPENDINGSTATUS[50]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS51 (CFGINTERRUPTMSIPENDINGSTATUS_IN[51], CFGINTERRUPTMSIPENDINGSTATUS[51]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS52 (CFGINTERRUPTMSIPENDINGSTATUS_IN[52], CFGINTERRUPTMSIPENDINGSTATUS[52]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS53 (CFGINTERRUPTMSIPENDINGSTATUS_IN[53], CFGINTERRUPTMSIPENDINGSTATUS[53]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS54 (CFGINTERRUPTMSIPENDINGSTATUS_IN[54], CFGINTERRUPTMSIPENDINGSTATUS[54]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS55 (CFGINTERRUPTMSIPENDINGSTATUS_IN[55], CFGINTERRUPTMSIPENDINGSTATUS[55]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS56 (CFGINTERRUPTMSIPENDINGSTATUS_IN[56], CFGINTERRUPTMSIPENDINGSTATUS[56]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS57 (CFGINTERRUPTMSIPENDINGSTATUS_IN[57], CFGINTERRUPTMSIPENDINGSTATUS[57]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS58 (CFGINTERRUPTMSIPENDINGSTATUS_IN[58], CFGINTERRUPTMSIPENDINGSTATUS[58]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS59 (CFGINTERRUPTMSIPENDINGSTATUS_IN[59], CFGINTERRUPTMSIPENDINGSTATUS[59]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS6 (CFGINTERRUPTMSIPENDINGSTATUS_IN[6], CFGINTERRUPTMSIPENDINGSTATUS[6]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS60 (CFGINTERRUPTMSIPENDINGSTATUS_IN[60], CFGINTERRUPTMSIPENDINGSTATUS[60]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS61 (CFGINTERRUPTMSIPENDINGSTATUS_IN[61], CFGINTERRUPTMSIPENDINGSTATUS[61]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS62 (CFGINTERRUPTMSIPENDINGSTATUS_IN[62], CFGINTERRUPTMSIPENDINGSTATUS[62]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS63 (CFGINTERRUPTMSIPENDINGSTATUS_IN[63], CFGINTERRUPTMSIPENDINGSTATUS[63]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS7 (CFGINTERRUPTMSIPENDINGSTATUS_IN[7], CFGINTERRUPTMSIPENDINGSTATUS[7]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS8 (CFGINTERRUPTMSIPENDINGSTATUS_IN[8], CFGINTERRUPTMSIPENDINGSTATUS[8]);
  buf B_CFGINTERRUPTMSIPENDINGSTATUS9 (CFGINTERRUPTMSIPENDINGSTATUS_IN[9], CFGINTERRUPTMSIPENDINGSTATUS[9]);
  buf B_CFGINTERRUPTMSISELECT0 (CFGINTERRUPTMSISELECT_IN[0], CFGINTERRUPTMSISELECT[0]);
  buf B_CFGINTERRUPTMSISELECT1 (CFGINTERRUPTMSISELECT_IN[1], CFGINTERRUPTMSISELECT[1]);
  buf B_CFGINTERRUPTMSISELECT2 (CFGINTERRUPTMSISELECT_IN[2], CFGINTERRUPTMSISELECT[2]);
  buf B_CFGINTERRUPTMSISELECT3 (CFGINTERRUPTMSISELECT_IN[3], CFGINTERRUPTMSISELECT[3]);
  buf B_CFGINTERRUPTMSITPHPRESENT (CFGINTERRUPTMSITPHPRESENT_IN, CFGINTERRUPTMSITPHPRESENT);
  buf B_CFGINTERRUPTMSITPHSTTAG0 (CFGINTERRUPTMSITPHSTTAG_IN[0], CFGINTERRUPTMSITPHSTTAG[0]);
  buf B_CFGINTERRUPTMSITPHSTTAG1 (CFGINTERRUPTMSITPHSTTAG_IN[1], CFGINTERRUPTMSITPHSTTAG[1]);
  buf B_CFGINTERRUPTMSITPHSTTAG2 (CFGINTERRUPTMSITPHSTTAG_IN[2], CFGINTERRUPTMSITPHSTTAG[2]);
  buf B_CFGINTERRUPTMSITPHSTTAG3 (CFGINTERRUPTMSITPHSTTAG_IN[3], CFGINTERRUPTMSITPHSTTAG[3]);
  buf B_CFGINTERRUPTMSITPHSTTAG4 (CFGINTERRUPTMSITPHSTTAG_IN[4], CFGINTERRUPTMSITPHSTTAG[4]);
  buf B_CFGINTERRUPTMSITPHSTTAG5 (CFGINTERRUPTMSITPHSTTAG_IN[5], CFGINTERRUPTMSITPHSTTAG[5]);
  buf B_CFGINTERRUPTMSITPHSTTAG6 (CFGINTERRUPTMSITPHSTTAG_IN[6], CFGINTERRUPTMSITPHSTTAG[6]);
  buf B_CFGINTERRUPTMSITPHSTTAG7 (CFGINTERRUPTMSITPHSTTAG_IN[7], CFGINTERRUPTMSITPHSTTAG[7]);
  buf B_CFGINTERRUPTMSITPHSTTAG8 (CFGINTERRUPTMSITPHSTTAG_IN[8], CFGINTERRUPTMSITPHSTTAG[8]);
  buf B_CFGINTERRUPTMSITPHTYPE0 (CFGINTERRUPTMSITPHTYPE_IN[0], CFGINTERRUPTMSITPHTYPE[0]);
  buf B_CFGINTERRUPTMSITPHTYPE1 (CFGINTERRUPTMSITPHTYPE_IN[1], CFGINTERRUPTMSITPHTYPE[1]);
  buf B_CFGINTERRUPTMSIXADDRESS0 (CFGINTERRUPTMSIXADDRESS_IN[0], CFGINTERRUPTMSIXADDRESS[0]);
  buf B_CFGINTERRUPTMSIXADDRESS1 (CFGINTERRUPTMSIXADDRESS_IN[1], CFGINTERRUPTMSIXADDRESS[1]);
  buf B_CFGINTERRUPTMSIXADDRESS10 (CFGINTERRUPTMSIXADDRESS_IN[10], CFGINTERRUPTMSIXADDRESS[10]);
  buf B_CFGINTERRUPTMSIXADDRESS11 (CFGINTERRUPTMSIXADDRESS_IN[11], CFGINTERRUPTMSIXADDRESS[11]);
  buf B_CFGINTERRUPTMSIXADDRESS12 (CFGINTERRUPTMSIXADDRESS_IN[12], CFGINTERRUPTMSIXADDRESS[12]);
  buf B_CFGINTERRUPTMSIXADDRESS13 (CFGINTERRUPTMSIXADDRESS_IN[13], CFGINTERRUPTMSIXADDRESS[13]);
  buf B_CFGINTERRUPTMSIXADDRESS14 (CFGINTERRUPTMSIXADDRESS_IN[14], CFGINTERRUPTMSIXADDRESS[14]);
  buf B_CFGINTERRUPTMSIXADDRESS15 (CFGINTERRUPTMSIXADDRESS_IN[15], CFGINTERRUPTMSIXADDRESS[15]);
  buf B_CFGINTERRUPTMSIXADDRESS16 (CFGINTERRUPTMSIXADDRESS_IN[16], CFGINTERRUPTMSIXADDRESS[16]);
  buf B_CFGINTERRUPTMSIXADDRESS17 (CFGINTERRUPTMSIXADDRESS_IN[17], CFGINTERRUPTMSIXADDRESS[17]);
  buf B_CFGINTERRUPTMSIXADDRESS18 (CFGINTERRUPTMSIXADDRESS_IN[18], CFGINTERRUPTMSIXADDRESS[18]);
  buf B_CFGINTERRUPTMSIXADDRESS19 (CFGINTERRUPTMSIXADDRESS_IN[19], CFGINTERRUPTMSIXADDRESS[19]);
  buf B_CFGINTERRUPTMSIXADDRESS2 (CFGINTERRUPTMSIXADDRESS_IN[2], CFGINTERRUPTMSIXADDRESS[2]);
  buf B_CFGINTERRUPTMSIXADDRESS20 (CFGINTERRUPTMSIXADDRESS_IN[20], CFGINTERRUPTMSIXADDRESS[20]);
  buf B_CFGINTERRUPTMSIXADDRESS21 (CFGINTERRUPTMSIXADDRESS_IN[21], CFGINTERRUPTMSIXADDRESS[21]);
  buf B_CFGINTERRUPTMSIXADDRESS22 (CFGINTERRUPTMSIXADDRESS_IN[22], CFGINTERRUPTMSIXADDRESS[22]);
  buf B_CFGINTERRUPTMSIXADDRESS23 (CFGINTERRUPTMSIXADDRESS_IN[23], CFGINTERRUPTMSIXADDRESS[23]);
  buf B_CFGINTERRUPTMSIXADDRESS24 (CFGINTERRUPTMSIXADDRESS_IN[24], CFGINTERRUPTMSIXADDRESS[24]);
  buf B_CFGINTERRUPTMSIXADDRESS25 (CFGINTERRUPTMSIXADDRESS_IN[25], CFGINTERRUPTMSIXADDRESS[25]);
  buf B_CFGINTERRUPTMSIXADDRESS26 (CFGINTERRUPTMSIXADDRESS_IN[26], CFGINTERRUPTMSIXADDRESS[26]);
  buf B_CFGINTERRUPTMSIXADDRESS27 (CFGINTERRUPTMSIXADDRESS_IN[27], CFGINTERRUPTMSIXADDRESS[27]);
  buf B_CFGINTERRUPTMSIXADDRESS28 (CFGINTERRUPTMSIXADDRESS_IN[28], CFGINTERRUPTMSIXADDRESS[28]);
  buf B_CFGINTERRUPTMSIXADDRESS29 (CFGINTERRUPTMSIXADDRESS_IN[29], CFGINTERRUPTMSIXADDRESS[29]);
  buf B_CFGINTERRUPTMSIXADDRESS3 (CFGINTERRUPTMSIXADDRESS_IN[3], CFGINTERRUPTMSIXADDRESS[3]);
  buf B_CFGINTERRUPTMSIXADDRESS30 (CFGINTERRUPTMSIXADDRESS_IN[30], CFGINTERRUPTMSIXADDRESS[30]);
  buf B_CFGINTERRUPTMSIXADDRESS31 (CFGINTERRUPTMSIXADDRESS_IN[31], CFGINTERRUPTMSIXADDRESS[31]);
  buf B_CFGINTERRUPTMSIXADDRESS32 (CFGINTERRUPTMSIXADDRESS_IN[32], CFGINTERRUPTMSIXADDRESS[32]);
  buf B_CFGINTERRUPTMSIXADDRESS33 (CFGINTERRUPTMSIXADDRESS_IN[33], CFGINTERRUPTMSIXADDRESS[33]);
  buf B_CFGINTERRUPTMSIXADDRESS34 (CFGINTERRUPTMSIXADDRESS_IN[34], CFGINTERRUPTMSIXADDRESS[34]);
  buf B_CFGINTERRUPTMSIXADDRESS35 (CFGINTERRUPTMSIXADDRESS_IN[35], CFGINTERRUPTMSIXADDRESS[35]);
  buf B_CFGINTERRUPTMSIXADDRESS36 (CFGINTERRUPTMSIXADDRESS_IN[36], CFGINTERRUPTMSIXADDRESS[36]);
  buf B_CFGINTERRUPTMSIXADDRESS37 (CFGINTERRUPTMSIXADDRESS_IN[37], CFGINTERRUPTMSIXADDRESS[37]);
  buf B_CFGINTERRUPTMSIXADDRESS38 (CFGINTERRUPTMSIXADDRESS_IN[38], CFGINTERRUPTMSIXADDRESS[38]);
  buf B_CFGINTERRUPTMSIXADDRESS39 (CFGINTERRUPTMSIXADDRESS_IN[39], CFGINTERRUPTMSIXADDRESS[39]);
  buf B_CFGINTERRUPTMSIXADDRESS4 (CFGINTERRUPTMSIXADDRESS_IN[4], CFGINTERRUPTMSIXADDRESS[4]);
  buf B_CFGINTERRUPTMSIXADDRESS40 (CFGINTERRUPTMSIXADDRESS_IN[40], CFGINTERRUPTMSIXADDRESS[40]);
  buf B_CFGINTERRUPTMSIXADDRESS41 (CFGINTERRUPTMSIXADDRESS_IN[41], CFGINTERRUPTMSIXADDRESS[41]);
  buf B_CFGINTERRUPTMSIXADDRESS42 (CFGINTERRUPTMSIXADDRESS_IN[42], CFGINTERRUPTMSIXADDRESS[42]);
  buf B_CFGINTERRUPTMSIXADDRESS43 (CFGINTERRUPTMSIXADDRESS_IN[43], CFGINTERRUPTMSIXADDRESS[43]);
  buf B_CFGINTERRUPTMSIXADDRESS44 (CFGINTERRUPTMSIXADDRESS_IN[44], CFGINTERRUPTMSIXADDRESS[44]);
  buf B_CFGINTERRUPTMSIXADDRESS45 (CFGINTERRUPTMSIXADDRESS_IN[45], CFGINTERRUPTMSIXADDRESS[45]);
  buf B_CFGINTERRUPTMSIXADDRESS46 (CFGINTERRUPTMSIXADDRESS_IN[46], CFGINTERRUPTMSIXADDRESS[46]);
  buf B_CFGINTERRUPTMSIXADDRESS47 (CFGINTERRUPTMSIXADDRESS_IN[47], CFGINTERRUPTMSIXADDRESS[47]);
  buf B_CFGINTERRUPTMSIXADDRESS48 (CFGINTERRUPTMSIXADDRESS_IN[48], CFGINTERRUPTMSIXADDRESS[48]);
  buf B_CFGINTERRUPTMSIXADDRESS49 (CFGINTERRUPTMSIXADDRESS_IN[49], CFGINTERRUPTMSIXADDRESS[49]);
  buf B_CFGINTERRUPTMSIXADDRESS5 (CFGINTERRUPTMSIXADDRESS_IN[5], CFGINTERRUPTMSIXADDRESS[5]);
  buf B_CFGINTERRUPTMSIXADDRESS50 (CFGINTERRUPTMSIXADDRESS_IN[50], CFGINTERRUPTMSIXADDRESS[50]);
  buf B_CFGINTERRUPTMSIXADDRESS51 (CFGINTERRUPTMSIXADDRESS_IN[51], CFGINTERRUPTMSIXADDRESS[51]);
  buf B_CFGINTERRUPTMSIXADDRESS52 (CFGINTERRUPTMSIXADDRESS_IN[52], CFGINTERRUPTMSIXADDRESS[52]);
  buf B_CFGINTERRUPTMSIXADDRESS53 (CFGINTERRUPTMSIXADDRESS_IN[53], CFGINTERRUPTMSIXADDRESS[53]);
  buf B_CFGINTERRUPTMSIXADDRESS54 (CFGINTERRUPTMSIXADDRESS_IN[54], CFGINTERRUPTMSIXADDRESS[54]);
  buf B_CFGINTERRUPTMSIXADDRESS55 (CFGINTERRUPTMSIXADDRESS_IN[55], CFGINTERRUPTMSIXADDRESS[55]);
  buf B_CFGINTERRUPTMSIXADDRESS56 (CFGINTERRUPTMSIXADDRESS_IN[56], CFGINTERRUPTMSIXADDRESS[56]);
  buf B_CFGINTERRUPTMSIXADDRESS57 (CFGINTERRUPTMSIXADDRESS_IN[57], CFGINTERRUPTMSIXADDRESS[57]);
  buf B_CFGINTERRUPTMSIXADDRESS58 (CFGINTERRUPTMSIXADDRESS_IN[58], CFGINTERRUPTMSIXADDRESS[58]);
  buf B_CFGINTERRUPTMSIXADDRESS59 (CFGINTERRUPTMSIXADDRESS_IN[59], CFGINTERRUPTMSIXADDRESS[59]);
  buf B_CFGINTERRUPTMSIXADDRESS6 (CFGINTERRUPTMSIXADDRESS_IN[6], CFGINTERRUPTMSIXADDRESS[6]);
  buf B_CFGINTERRUPTMSIXADDRESS60 (CFGINTERRUPTMSIXADDRESS_IN[60], CFGINTERRUPTMSIXADDRESS[60]);
  buf B_CFGINTERRUPTMSIXADDRESS61 (CFGINTERRUPTMSIXADDRESS_IN[61], CFGINTERRUPTMSIXADDRESS[61]);
  buf B_CFGINTERRUPTMSIXADDRESS62 (CFGINTERRUPTMSIXADDRESS_IN[62], CFGINTERRUPTMSIXADDRESS[62]);
  buf B_CFGINTERRUPTMSIXADDRESS63 (CFGINTERRUPTMSIXADDRESS_IN[63], CFGINTERRUPTMSIXADDRESS[63]);
  buf B_CFGINTERRUPTMSIXADDRESS7 (CFGINTERRUPTMSIXADDRESS_IN[7], CFGINTERRUPTMSIXADDRESS[7]);
  buf B_CFGINTERRUPTMSIXADDRESS8 (CFGINTERRUPTMSIXADDRESS_IN[8], CFGINTERRUPTMSIXADDRESS[8]);
  buf B_CFGINTERRUPTMSIXADDRESS9 (CFGINTERRUPTMSIXADDRESS_IN[9], CFGINTERRUPTMSIXADDRESS[9]);
  buf B_CFGINTERRUPTMSIXDATA0 (CFGINTERRUPTMSIXDATA_IN[0], CFGINTERRUPTMSIXDATA[0]);
  buf B_CFGINTERRUPTMSIXDATA1 (CFGINTERRUPTMSIXDATA_IN[1], CFGINTERRUPTMSIXDATA[1]);
  buf B_CFGINTERRUPTMSIXDATA10 (CFGINTERRUPTMSIXDATA_IN[10], CFGINTERRUPTMSIXDATA[10]);
  buf B_CFGINTERRUPTMSIXDATA11 (CFGINTERRUPTMSIXDATA_IN[11], CFGINTERRUPTMSIXDATA[11]);
  buf B_CFGINTERRUPTMSIXDATA12 (CFGINTERRUPTMSIXDATA_IN[12], CFGINTERRUPTMSIXDATA[12]);
  buf B_CFGINTERRUPTMSIXDATA13 (CFGINTERRUPTMSIXDATA_IN[13], CFGINTERRUPTMSIXDATA[13]);
  buf B_CFGINTERRUPTMSIXDATA14 (CFGINTERRUPTMSIXDATA_IN[14], CFGINTERRUPTMSIXDATA[14]);
  buf B_CFGINTERRUPTMSIXDATA15 (CFGINTERRUPTMSIXDATA_IN[15], CFGINTERRUPTMSIXDATA[15]);
  buf B_CFGINTERRUPTMSIXDATA16 (CFGINTERRUPTMSIXDATA_IN[16], CFGINTERRUPTMSIXDATA[16]);
  buf B_CFGINTERRUPTMSIXDATA17 (CFGINTERRUPTMSIXDATA_IN[17], CFGINTERRUPTMSIXDATA[17]);
  buf B_CFGINTERRUPTMSIXDATA18 (CFGINTERRUPTMSIXDATA_IN[18], CFGINTERRUPTMSIXDATA[18]);
  buf B_CFGINTERRUPTMSIXDATA19 (CFGINTERRUPTMSIXDATA_IN[19], CFGINTERRUPTMSIXDATA[19]);
  buf B_CFGINTERRUPTMSIXDATA2 (CFGINTERRUPTMSIXDATA_IN[2], CFGINTERRUPTMSIXDATA[2]);
  buf B_CFGINTERRUPTMSIXDATA20 (CFGINTERRUPTMSIXDATA_IN[20], CFGINTERRUPTMSIXDATA[20]);
  buf B_CFGINTERRUPTMSIXDATA21 (CFGINTERRUPTMSIXDATA_IN[21], CFGINTERRUPTMSIXDATA[21]);
  buf B_CFGINTERRUPTMSIXDATA22 (CFGINTERRUPTMSIXDATA_IN[22], CFGINTERRUPTMSIXDATA[22]);
  buf B_CFGINTERRUPTMSIXDATA23 (CFGINTERRUPTMSIXDATA_IN[23], CFGINTERRUPTMSIXDATA[23]);
  buf B_CFGINTERRUPTMSIXDATA24 (CFGINTERRUPTMSIXDATA_IN[24], CFGINTERRUPTMSIXDATA[24]);
  buf B_CFGINTERRUPTMSIXDATA25 (CFGINTERRUPTMSIXDATA_IN[25], CFGINTERRUPTMSIXDATA[25]);
  buf B_CFGINTERRUPTMSIXDATA26 (CFGINTERRUPTMSIXDATA_IN[26], CFGINTERRUPTMSIXDATA[26]);
  buf B_CFGINTERRUPTMSIXDATA27 (CFGINTERRUPTMSIXDATA_IN[27], CFGINTERRUPTMSIXDATA[27]);
  buf B_CFGINTERRUPTMSIXDATA28 (CFGINTERRUPTMSIXDATA_IN[28], CFGINTERRUPTMSIXDATA[28]);
  buf B_CFGINTERRUPTMSIXDATA29 (CFGINTERRUPTMSIXDATA_IN[29], CFGINTERRUPTMSIXDATA[29]);
  buf B_CFGINTERRUPTMSIXDATA3 (CFGINTERRUPTMSIXDATA_IN[3], CFGINTERRUPTMSIXDATA[3]);
  buf B_CFGINTERRUPTMSIXDATA30 (CFGINTERRUPTMSIXDATA_IN[30], CFGINTERRUPTMSIXDATA[30]);
  buf B_CFGINTERRUPTMSIXDATA31 (CFGINTERRUPTMSIXDATA_IN[31], CFGINTERRUPTMSIXDATA[31]);
  buf B_CFGINTERRUPTMSIXDATA4 (CFGINTERRUPTMSIXDATA_IN[4], CFGINTERRUPTMSIXDATA[4]);
  buf B_CFGINTERRUPTMSIXDATA5 (CFGINTERRUPTMSIXDATA_IN[5], CFGINTERRUPTMSIXDATA[5]);
  buf B_CFGINTERRUPTMSIXDATA6 (CFGINTERRUPTMSIXDATA_IN[6], CFGINTERRUPTMSIXDATA[6]);
  buf B_CFGINTERRUPTMSIXDATA7 (CFGINTERRUPTMSIXDATA_IN[7], CFGINTERRUPTMSIXDATA[7]);
  buf B_CFGINTERRUPTMSIXDATA8 (CFGINTERRUPTMSIXDATA_IN[8], CFGINTERRUPTMSIXDATA[8]);
  buf B_CFGINTERRUPTMSIXDATA9 (CFGINTERRUPTMSIXDATA_IN[9], CFGINTERRUPTMSIXDATA[9]);
  buf B_CFGINTERRUPTMSIXINT (CFGINTERRUPTMSIXINT_IN, CFGINTERRUPTMSIXINT);
  buf B_CFGINTERRUPTPENDING0 (CFGINTERRUPTPENDING_IN[0], CFGINTERRUPTPENDING[0]);
  buf B_CFGINTERRUPTPENDING1 (CFGINTERRUPTPENDING_IN[1], CFGINTERRUPTPENDING[1]);
  buf B_CFGLINKTRAININGENABLE (CFGLINKTRAININGENABLE_IN, CFGLINKTRAININGENABLE);
  buf B_CFGMCUPDATEREQUEST (CFGMCUPDATEREQUEST_IN, CFGMCUPDATEREQUEST);
  buf B_CFGMGMTADDR0 (CFGMGMTADDR_IN[0], CFGMGMTADDR[0]);
  buf B_CFGMGMTADDR1 (CFGMGMTADDR_IN[1], CFGMGMTADDR[1]);
  buf B_CFGMGMTADDR10 (CFGMGMTADDR_IN[10], CFGMGMTADDR[10]);
  buf B_CFGMGMTADDR11 (CFGMGMTADDR_IN[11], CFGMGMTADDR[11]);
  buf B_CFGMGMTADDR12 (CFGMGMTADDR_IN[12], CFGMGMTADDR[12]);
  buf B_CFGMGMTADDR13 (CFGMGMTADDR_IN[13], CFGMGMTADDR[13]);
  buf B_CFGMGMTADDR14 (CFGMGMTADDR_IN[14], CFGMGMTADDR[14]);
  buf B_CFGMGMTADDR15 (CFGMGMTADDR_IN[15], CFGMGMTADDR[15]);
  buf B_CFGMGMTADDR16 (CFGMGMTADDR_IN[16], CFGMGMTADDR[16]);
  buf B_CFGMGMTADDR17 (CFGMGMTADDR_IN[17], CFGMGMTADDR[17]);
  buf B_CFGMGMTADDR18 (CFGMGMTADDR_IN[18], CFGMGMTADDR[18]);
  buf B_CFGMGMTADDR2 (CFGMGMTADDR_IN[2], CFGMGMTADDR[2]);
  buf B_CFGMGMTADDR3 (CFGMGMTADDR_IN[3], CFGMGMTADDR[3]);
  buf B_CFGMGMTADDR4 (CFGMGMTADDR_IN[4], CFGMGMTADDR[4]);
  buf B_CFGMGMTADDR5 (CFGMGMTADDR_IN[5], CFGMGMTADDR[5]);
  buf B_CFGMGMTADDR6 (CFGMGMTADDR_IN[6], CFGMGMTADDR[6]);
  buf B_CFGMGMTADDR7 (CFGMGMTADDR_IN[7], CFGMGMTADDR[7]);
  buf B_CFGMGMTADDR8 (CFGMGMTADDR_IN[8], CFGMGMTADDR[8]);
  buf B_CFGMGMTADDR9 (CFGMGMTADDR_IN[9], CFGMGMTADDR[9]);
  buf B_CFGMGMTBYTEENABLE0 (CFGMGMTBYTEENABLE_IN[0], CFGMGMTBYTEENABLE[0]);
  buf B_CFGMGMTBYTEENABLE1 (CFGMGMTBYTEENABLE_IN[1], CFGMGMTBYTEENABLE[1]);
  buf B_CFGMGMTBYTEENABLE2 (CFGMGMTBYTEENABLE_IN[2], CFGMGMTBYTEENABLE[2]);
  buf B_CFGMGMTBYTEENABLE3 (CFGMGMTBYTEENABLE_IN[3], CFGMGMTBYTEENABLE[3]);
  buf B_CFGMGMTREAD (CFGMGMTREAD_IN, CFGMGMTREAD);
  buf B_CFGMGMTTYPE1CFGREGACCESS (CFGMGMTTYPE1CFGREGACCESS_IN, CFGMGMTTYPE1CFGREGACCESS);
  buf B_CFGMGMTWRITE (CFGMGMTWRITE_IN, CFGMGMTWRITE);
  buf B_CFGMGMTWRITEDATA0 (CFGMGMTWRITEDATA_IN[0], CFGMGMTWRITEDATA[0]);
  buf B_CFGMGMTWRITEDATA1 (CFGMGMTWRITEDATA_IN[1], CFGMGMTWRITEDATA[1]);
  buf B_CFGMGMTWRITEDATA10 (CFGMGMTWRITEDATA_IN[10], CFGMGMTWRITEDATA[10]);
  buf B_CFGMGMTWRITEDATA11 (CFGMGMTWRITEDATA_IN[11], CFGMGMTWRITEDATA[11]);
  buf B_CFGMGMTWRITEDATA12 (CFGMGMTWRITEDATA_IN[12], CFGMGMTWRITEDATA[12]);
  buf B_CFGMGMTWRITEDATA13 (CFGMGMTWRITEDATA_IN[13], CFGMGMTWRITEDATA[13]);
  buf B_CFGMGMTWRITEDATA14 (CFGMGMTWRITEDATA_IN[14], CFGMGMTWRITEDATA[14]);
  buf B_CFGMGMTWRITEDATA15 (CFGMGMTWRITEDATA_IN[15], CFGMGMTWRITEDATA[15]);
  buf B_CFGMGMTWRITEDATA16 (CFGMGMTWRITEDATA_IN[16], CFGMGMTWRITEDATA[16]);
  buf B_CFGMGMTWRITEDATA17 (CFGMGMTWRITEDATA_IN[17], CFGMGMTWRITEDATA[17]);
  buf B_CFGMGMTWRITEDATA18 (CFGMGMTWRITEDATA_IN[18], CFGMGMTWRITEDATA[18]);
  buf B_CFGMGMTWRITEDATA19 (CFGMGMTWRITEDATA_IN[19], CFGMGMTWRITEDATA[19]);
  buf B_CFGMGMTWRITEDATA2 (CFGMGMTWRITEDATA_IN[2], CFGMGMTWRITEDATA[2]);
  buf B_CFGMGMTWRITEDATA20 (CFGMGMTWRITEDATA_IN[20], CFGMGMTWRITEDATA[20]);
  buf B_CFGMGMTWRITEDATA21 (CFGMGMTWRITEDATA_IN[21], CFGMGMTWRITEDATA[21]);
  buf B_CFGMGMTWRITEDATA22 (CFGMGMTWRITEDATA_IN[22], CFGMGMTWRITEDATA[22]);
  buf B_CFGMGMTWRITEDATA23 (CFGMGMTWRITEDATA_IN[23], CFGMGMTWRITEDATA[23]);
  buf B_CFGMGMTWRITEDATA24 (CFGMGMTWRITEDATA_IN[24], CFGMGMTWRITEDATA[24]);
  buf B_CFGMGMTWRITEDATA25 (CFGMGMTWRITEDATA_IN[25], CFGMGMTWRITEDATA[25]);
  buf B_CFGMGMTWRITEDATA26 (CFGMGMTWRITEDATA_IN[26], CFGMGMTWRITEDATA[26]);
  buf B_CFGMGMTWRITEDATA27 (CFGMGMTWRITEDATA_IN[27], CFGMGMTWRITEDATA[27]);
  buf B_CFGMGMTWRITEDATA28 (CFGMGMTWRITEDATA_IN[28], CFGMGMTWRITEDATA[28]);
  buf B_CFGMGMTWRITEDATA29 (CFGMGMTWRITEDATA_IN[29], CFGMGMTWRITEDATA[29]);
  buf B_CFGMGMTWRITEDATA3 (CFGMGMTWRITEDATA_IN[3], CFGMGMTWRITEDATA[3]);
  buf B_CFGMGMTWRITEDATA30 (CFGMGMTWRITEDATA_IN[30], CFGMGMTWRITEDATA[30]);
  buf B_CFGMGMTWRITEDATA31 (CFGMGMTWRITEDATA_IN[31], CFGMGMTWRITEDATA[31]);
  buf B_CFGMGMTWRITEDATA4 (CFGMGMTWRITEDATA_IN[4], CFGMGMTWRITEDATA[4]);
  buf B_CFGMGMTWRITEDATA5 (CFGMGMTWRITEDATA_IN[5], CFGMGMTWRITEDATA[5]);
  buf B_CFGMGMTWRITEDATA6 (CFGMGMTWRITEDATA_IN[6], CFGMGMTWRITEDATA[6]);
  buf B_CFGMGMTWRITEDATA7 (CFGMGMTWRITEDATA_IN[7], CFGMGMTWRITEDATA[7]);
  buf B_CFGMGMTWRITEDATA8 (CFGMGMTWRITEDATA_IN[8], CFGMGMTWRITEDATA[8]);
  buf B_CFGMGMTWRITEDATA9 (CFGMGMTWRITEDATA_IN[9], CFGMGMTWRITEDATA[9]);
  buf B_CFGMSGTRANSMIT (CFGMSGTRANSMIT_IN, CFGMSGTRANSMIT);
  buf B_CFGMSGTRANSMITDATA0 (CFGMSGTRANSMITDATA_IN[0], CFGMSGTRANSMITDATA[0]);
  buf B_CFGMSGTRANSMITDATA1 (CFGMSGTRANSMITDATA_IN[1], CFGMSGTRANSMITDATA[1]);
  buf B_CFGMSGTRANSMITDATA10 (CFGMSGTRANSMITDATA_IN[10], CFGMSGTRANSMITDATA[10]);
  buf B_CFGMSGTRANSMITDATA11 (CFGMSGTRANSMITDATA_IN[11], CFGMSGTRANSMITDATA[11]);
  buf B_CFGMSGTRANSMITDATA12 (CFGMSGTRANSMITDATA_IN[12], CFGMSGTRANSMITDATA[12]);
  buf B_CFGMSGTRANSMITDATA13 (CFGMSGTRANSMITDATA_IN[13], CFGMSGTRANSMITDATA[13]);
  buf B_CFGMSGTRANSMITDATA14 (CFGMSGTRANSMITDATA_IN[14], CFGMSGTRANSMITDATA[14]);
  buf B_CFGMSGTRANSMITDATA15 (CFGMSGTRANSMITDATA_IN[15], CFGMSGTRANSMITDATA[15]);
  buf B_CFGMSGTRANSMITDATA16 (CFGMSGTRANSMITDATA_IN[16], CFGMSGTRANSMITDATA[16]);
  buf B_CFGMSGTRANSMITDATA17 (CFGMSGTRANSMITDATA_IN[17], CFGMSGTRANSMITDATA[17]);
  buf B_CFGMSGTRANSMITDATA18 (CFGMSGTRANSMITDATA_IN[18], CFGMSGTRANSMITDATA[18]);
  buf B_CFGMSGTRANSMITDATA19 (CFGMSGTRANSMITDATA_IN[19], CFGMSGTRANSMITDATA[19]);
  buf B_CFGMSGTRANSMITDATA2 (CFGMSGTRANSMITDATA_IN[2], CFGMSGTRANSMITDATA[2]);
  buf B_CFGMSGTRANSMITDATA20 (CFGMSGTRANSMITDATA_IN[20], CFGMSGTRANSMITDATA[20]);
  buf B_CFGMSGTRANSMITDATA21 (CFGMSGTRANSMITDATA_IN[21], CFGMSGTRANSMITDATA[21]);
  buf B_CFGMSGTRANSMITDATA22 (CFGMSGTRANSMITDATA_IN[22], CFGMSGTRANSMITDATA[22]);
  buf B_CFGMSGTRANSMITDATA23 (CFGMSGTRANSMITDATA_IN[23], CFGMSGTRANSMITDATA[23]);
  buf B_CFGMSGTRANSMITDATA24 (CFGMSGTRANSMITDATA_IN[24], CFGMSGTRANSMITDATA[24]);
  buf B_CFGMSGTRANSMITDATA25 (CFGMSGTRANSMITDATA_IN[25], CFGMSGTRANSMITDATA[25]);
  buf B_CFGMSGTRANSMITDATA26 (CFGMSGTRANSMITDATA_IN[26], CFGMSGTRANSMITDATA[26]);
  buf B_CFGMSGTRANSMITDATA27 (CFGMSGTRANSMITDATA_IN[27], CFGMSGTRANSMITDATA[27]);
  buf B_CFGMSGTRANSMITDATA28 (CFGMSGTRANSMITDATA_IN[28], CFGMSGTRANSMITDATA[28]);
  buf B_CFGMSGTRANSMITDATA29 (CFGMSGTRANSMITDATA_IN[29], CFGMSGTRANSMITDATA[29]);
  buf B_CFGMSGTRANSMITDATA3 (CFGMSGTRANSMITDATA_IN[3], CFGMSGTRANSMITDATA[3]);
  buf B_CFGMSGTRANSMITDATA30 (CFGMSGTRANSMITDATA_IN[30], CFGMSGTRANSMITDATA[30]);
  buf B_CFGMSGTRANSMITDATA31 (CFGMSGTRANSMITDATA_IN[31], CFGMSGTRANSMITDATA[31]);
  buf B_CFGMSGTRANSMITDATA4 (CFGMSGTRANSMITDATA_IN[4], CFGMSGTRANSMITDATA[4]);
  buf B_CFGMSGTRANSMITDATA5 (CFGMSGTRANSMITDATA_IN[5], CFGMSGTRANSMITDATA[5]);
  buf B_CFGMSGTRANSMITDATA6 (CFGMSGTRANSMITDATA_IN[6], CFGMSGTRANSMITDATA[6]);
  buf B_CFGMSGTRANSMITDATA7 (CFGMSGTRANSMITDATA_IN[7], CFGMSGTRANSMITDATA[7]);
  buf B_CFGMSGTRANSMITDATA8 (CFGMSGTRANSMITDATA_IN[8], CFGMSGTRANSMITDATA[8]);
  buf B_CFGMSGTRANSMITDATA9 (CFGMSGTRANSMITDATA_IN[9], CFGMSGTRANSMITDATA[9]);
  buf B_CFGMSGTRANSMITTYPE0 (CFGMSGTRANSMITTYPE_IN[0], CFGMSGTRANSMITTYPE[0]);
  buf B_CFGMSGTRANSMITTYPE1 (CFGMSGTRANSMITTYPE_IN[1], CFGMSGTRANSMITTYPE[1]);
  buf B_CFGMSGTRANSMITTYPE2 (CFGMSGTRANSMITTYPE_IN[2], CFGMSGTRANSMITTYPE[2]);
  buf B_CFGPERFUNCSTATUSCONTROL0 (CFGPERFUNCSTATUSCONTROL_IN[0], CFGPERFUNCSTATUSCONTROL[0]);
  buf B_CFGPERFUNCSTATUSCONTROL1 (CFGPERFUNCSTATUSCONTROL_IN[1], CFGPERFUNCSTATUSCONTROL[1]);
  buf B_CFGPERFUNCSTATUSCONTROL2 (CFGPERFUNCSTATUSCONTROL_IN[2], CFGPERFUNCSTATUSCONTROL[2]);
  buf B_CFGPERFUNCTIONNUMBER0 (CFGPERFUNCTIONNUMBER_IN[0], CFGPERFUNCTIONNUMBER[0]);
  buf B_CFGPERFUNCTIONNUMBER1 (CFGPERFUNCTIONNUMBER_IN[1], CFGPERFUNCTIONNUMBER[1]);
  buf B_CFGPERFUNCTIONNUMBER2 (CFGPERFUNCTIONNUMBER_IN[2], CFGPERFUNCTIONNUMBER[2]);
  buf B_CFGPERFUNCTIONOUTPUTREQUEST (CFGPERFUNCTIONOUTPUTREQUEST_IN, CFGPERFUNCTIONOUTPUTREQUEST);
  buf B_CFGPOWERSTATECHANGEACK (CFGPOWERSTATECHANGEACK_IN, CFGPOWERSTATECHANGEACK);
  buf B_CFGREQPMTRANSITIONL23READY (CFGREQPMTRANSITIONL23READY_IN, CFGREQPMTRANSITIONL23READY);
  buf B_CFGREVID0 (CFGREVID_IN[0], CFGREVID[0]);
  buf B_CFGREVID1 (CFGREVID_IN[1], CFGREVID[1]);
  buf B_CFGREVID2 (CFGREVID_IN[2], CFGREVID[2]);
  buf B_CFGREVID3 (CFGREVID_IN[3], CFGREVID[3]);
  buf B_CFGREVID4 (CFGREVID_IN[4], CFGREVID[4]);
  buf B_CFGREVID5 (CFGREVID_IN[5], CFGREVID[5]);
  buf B_CFGREVID6 (CFGREVID_IN[6], CFGREVID[6]);
  buf B_CFGREVID7 (CFGREVID_IN[7], CFGREVID[7]);
  buf B_CFGSUBSYSID0 (CFGSUBSYSID_IN[0], CFGSUBSYSID[0]);
  buf B_CFGSUBSYSID1 (CFGSUBSYSID_IN[1], CFGSUBSYSID[1]);
  buf B_CFGSUBSYSID10 (CFGSUBSYSID_IN[10], CFGSUBSYSID[10]);
  buf B_CFGSUBSYSID11 (CFGSUBSYSID_IN[11], CFGSUBSYSID[11]);
  buf B_CFGSUBSYSID12 (CFGSUBSYSID_IN[12], CFGSUBSYSID[12]);
  buf B_CFGSUBSYSID13 (CFGSUBSYSID_IN[13], CFGSUBSYSID[13]);
  buf B_CFGSUBSYSID14 (CFGSUBSYSID_IN[14], CFGSUBSYSID[14]);
  buf B_CFGSUBSYSID15 (CFGSUBSYSID_IN[15], CFGSUBSYSID[15]);
  buf B_CFGSUBSYSID2 (CFGSUBSYSID_IN[2], CFGSUBSYSID[2]);
  buf B_CFGSUBSYSID3 (CFGSUBSYSID_IN[3], CFGSUBSYSID[3]);
  buf B_CFGSUBSYSID4 (CFGSUBSYSID_IN[4], CFGSUBSYSID[4]);
  buf B_CFGSUBSYSID5 (CFGSUBSYSID_IN[5], CFGSUBSYSID[5]);
  buf B_CFGSUBSYSID6 (CFGSUBSYSID_IN[6], CFGSUBSYSID[6]);
  buf B_CFGSUBSYSID7 (CFGSUBSYSID_IN[7], CFGSUBSYSID[7]);
  buf B_CFGSUBSYSID8 (CFGSUBSYSID_IN[8], CFGSUBSYSID[8]);
  buf B_CFGSUBSYSID9 (CFGSUBSYSID_IN[9], CFGSUBSYSID[9]);
  buf B_CFGSUBSYSVENDID0 (CFGSUBSYSVENDID_IN[0], CFGSUBSYSVENDID[0]);
  buf B_CFGSUBSYSVENDID1 (CFGSUBSYSVENDID_IN[1], CFGSUBSYSVENDID[1]);
  buf B_CFGSUBSYSVENDID10 (CFGSUBSYSVENDID_IN[10], CFGSUBSYSVENDID[10]);
  buf B_CFGSUBSYSVENDID11 (CFGSUBSYSVENDID_IN[11], CFGSUBSYSVENDID[11]);
  buf B_CFGSUBSYSVENDID12 (CFGSUBSYSVENDID_IN[12], CFGSUBSYSVENDID[12]);
  buf B_CFGSUBSYSVENDID13 (CFGSUBSYSVENDID_IN[13], CFGSUBSYSVENDID[13]);
  buf B_CFGSUBSYSVENDID14 (CFGSUBSYSVENDID_IN[14], CFGSUBSYSVENDID[14]);
  buf B_CFGSUBSYSVENDID15 (CFGSUBSYSVENDID_IN[15], CFGSUBSYSVENDID[15]);
  buf B_CFGSUBSYSVENDID2 (CFGSUBSYSVENDID_IN[2], CFGSUBSYSVENDID[2]);
  buf B_CFGSUBSYSVENDID3 (CFGSUBSYSVENDID_IN[3], CFGSUBSYSVENDID[3]);
  buf B_CFGSUBSYSVENDID4 (CFGSUBSYSVENDID_IN[4], CFGSUBSYSVENDID[4]);
  buf B_CFGSUBSYSVENDID5 (CFGSUBSYSVENDID_IN[5], CFGSUBSYSVENDID[5]);
  buf B_CFGSUBSYSVENDID6 (CFGSUBSYSVENDID_IN[6], CFGSUBSYSVENDID[6]);
  buf B_CFGSUBSYSVENDID7 (CFGSUBSYSVENDID_IN[7], CFGSUBSYSVENDID[7]);
  buf B_CFGSUBSYSVENDID8 (CFGSUBSYSVENDID_IN[8], CFGSUBSYSVENDID[8]);
  buf B_CFGSUBSYSVENDID9 (CFGSUBSYSVENDID_IN[9], CFGSUBSYSVENDID[9]);
  buf B_CFGTPHSTTREADDATA0 (CFGTPHSTTREADDATA_IN[0], CFGTPHSTTREADDATA[0]);
  buf B_CFGTPHSTTREADDATA1 (CFGTPHSTTREADDATA_IN[1], CFGTPHSTTREADDATA[1]);
  buf B_CFGTPHSTTREADDATA10 (CFGTPHSTTREADDATA_IN[10], CFGTPHSTTREADDATA[10]);
  buf B_CFGTPHSTTREADDATA11 (CFGTPHSTTREADDATA_IN[11], CFGTPHSTTREADDATA[11]);
  buf B_CFGTPHSTTREADDATA12 (CFGTPHSTTREADDATA_IN[12], CFGTPHSTTREADDATA[12]);
  buf B_CFGTPHSTTREADDATA13 (CFGTPHSTTREADDATA_IN[13], CFGTPHSTTREADDATA[13]);
  buf B_CFGTPHSTTREADDATA14 (CFGTPHSTTREADDATA_IN[14], CFGTPHSTTREADDATA[14]);
  buf B_CFGTPHSTTREADDATA15 (CFGTPHSTTREADDATA_IN[15], CFGTPHSTTREADDATA[15]);
  buf B_CFGTPHSTTREADDATA16 (CFGTPHSTTREADDATA_IN[16], CFGTPHSTTREADDATA[16]);
  buf B_CFGTPHSTTREADDATA17 (CFGTPHSTTREADDATA_IN[17], CFGTPHSTTREADDATA[17]);
  buf B_CFGTPHSTTREADDATA18 (CFGTPHSTTREADDATA_IN[18], CFGTPHSTTREADDATA[18]);
  buf B_CFGTPHSTTREADDATA19 (CFGTPHSTTREADDATA_IN[19], CFGTPHSTTREADDATA[19]);
  buf B_CFGTPHSTTREADDATA2 (CFGTPHSTTREADDATA_IN[2], CFGTPHSTTREADDATA[2]);
  buf B_CFGTPHSTTREADDATA20 (CFGTPHSTTREADDATA_IN[20], CFGTPHSTTREADDATA[20]);
  buf B_CFGTPHSTTREADDATA21 (CFGTPHSTTREADDATA_IN[21], CFGTPHSTTREADDATA[21]);
  buf B_CFGTPHSTTREADDATA22 (CFGTPHSTTREADDATA_IN[22], CFGTPHSTTREADDATA[22]);
  buf B_CFGTPHSTTREADDATA23 (CFGTPHSTTREADDATA_IN[23], CFGTPHSTTREADDATA[23]);
  buf B_CFGTPHSTTREADDATA24 (CFGTPHSTTREADDATA_IN[24], CFGTPHSTTREADDATA[24]);
  buf B_CFGTPHSTTREADDATA25 (CFGTPHSTTREADDATA_IN[25], CFGTPHSTTREADDATA[25]);
  buf B_CFGTPHSTTREADDATA26 (CFGTPHSTTREADDATA_IN[26], CFGTPHSTTREADDATA[26]);
  buf B_CFGTPHSTTREADDATA27 (CFGTPHSTTREADDATA_IN[27], CFGTPHSTTREADDATA[27]);
  buf B_CFGTPHSTTREADDATA28 (CFGTPHSTTREADDATA_IN[28], CFGTPHSTTREADDATA[28]);
  buf B_CFGTPHSTTREADDATA29 (CFGTPHSTTREADDATA_IN[29], CFGTPHSTTREADDATA[29]);
  buf B_CFGTPHSTTREADDATA3 (CFGTPHSTTREADDATA_IN[3], CFGTPHSTTREADDATA[3]);
  buf B_CFGTPHSTTREADDATA30 (CFGTPHSTTREADDATA_IN[30], CFGTPHSTTREADDATA[30]);
  buf B_CFGTPHSTTREADDATA31 (CFGTPHSTTREADDATA_IN[31], CFGTPHSTTREADDATA[31]);
  buf B_CFGTPHSTTREADDATA4 (CFGTPHSTTREADDATA_IN[4], CFGTPHSTTREADDATA[4]);
  buf B_CFGTPHSTTREADDATA5 (CFGTPHSTTREADDATA_IN[5], CFGTPHSTTREADDATA[5]);
  buf B_CFGTPHSTTREADDATA6 (CFGTPHSTTREADDATA_IN[6], CFGTPHSTTREADDATA[6]);
  buf B_CFGTPHSTTREADDATA7 (CFGTPHSTTREADDATA_IN[7], CFGTPHSTTREADDATA[7]);
  buf B_CFGTPHSTTREADDATA8 (CFGTPHSTTREADDATA_IN[8], CFGTPHSTTREADDATA[8]);
  buf B_CFGTPHSTTREADDATA9 (CFGTPHSTTREADDATA_IN[9], CFGTPHSTTREADDATA[9]);
  buf B_CFGTPHSTTREADDATAVALID (CFGTPHSTTREADDATAVALID_IN, CFGTPHSTTREADDATAVALID);
  buf B_CFGVENDID0 (CFGVENDID_IN[0], CFGVENDID[0]);
  buf B_CFGVENDID1 (CFGVENDID_IN[1], CFGVENDID[1]);
  buf B_CFGVENDID10 (CFGVENDID_IN[10], CFGVENDID[10]);
  buf B_CFGVENDID11 (CFGVENDID_IN[11], CFGVENDID[11]);
  buf B_CFGVENDID12 (CFGVENDID_IN[12], CFGVENDID[12]);
  buf B_CFGVENDID13 (CFGVENDID_IN[13], CFGVENDID[13]);
  buf B_CFGVENDID14 (CFGVENDID_IN[14], CFGVENDID[14]);
  buf B_CFGVENDID15 (CFGVENDID_IN[15], CFGVENDID[15]);
  buf B_CFGVENDID2 (CFGVENDID_IN[2], CFGVENDID[2]);
  buf B_CFGVENDID3 (CFGVENDID_IN[3], CFGVENDID[3]);
  buf B_CFGVENDID4 (CFGVENDID_IN[4], CFGVENDID[4]);
  buf B_CFGVENDID5 (CFGVENDID_IN[5], CFGVENDID[5]);
  buf B_CFGVENDID6 (CFGVENDID_IN[6], CFGVENDID[6]);
  buf B_CFGVENDID7 (CFGVENDID_IN[7], CFGVENDID[7]);
  buf B_CFGVENDID8 (CFGVENDID_IN[8], CFGVENDID[8]);
  buf B_CFGVENDID9 (CFGVENDID_IN[9], CFGVENDID[9]);
  buf B_CFGVFFLRDONE0 (CFGVFFLRDONE_IN[0], CFGVFFLRDONE[0]);
  buf B_CFGVFFLRDONE1 (CFGVFFLRDONE_IN[1], CFGVFFLRDONE[1]);
  buf B_CFGVFFLRDONE2 (CFGVFFLRDONE_IN[2], CFGVFFLRDONE[2]);
  buf B_CFGVFFLRDONE3 (CFGVFFLRDONE_IN[3], CFGVFFLRDONE[3]);
  buf B_CFGVFFLRDONE4 (CFGVFFLRDONE_IN[4], CFGVFFLRDONE[4]);
  buf B_CFGVFFLRDONE5 (CFGVFFLRDONE_IN[5], CFGVFFLRDONE[5]);
  buf B_CORECLK (CORECLK_IN, CORECLK);
  buf B_CORECLKMICOMPLETIONRAML (CORECLKMICOMPLETIONRAML_IN, CORECLKMICOMPLETIONRAML);
  buf B_CORECLKMICOMPLETIONRAMU (CORECLKMICOMPLETIONRAMU_IN, CORECLKMICOMPLETIONRAMU);
  buf B_CORECLKMIREPLAYRAM (CORECLKMIREPLAYRAM_IN, CORECLKMIREPLAYRAM);
  buf B_CORECLKMIREQUESTRAM (CORECLKMIREQUESTRAM_IN, CORECLKMIREQUESTRAM);
  buf B_DRPADDR0 (DRPADDR_IN[0], DRPADDR[0]);
  buf B_DRPADDR1 (DRPADDR_IN[1], DRPADDR[1]);
  buf B_DRPADDR10 (DRPADDR_IN[10], DRPADDR[10]);
  buf B_DRPADDR2 (DRPADDR_IN[2], DRPADDR[2]);
  buf B_DRPADDR3 (DRPADDR_IN[3], DRPADDR[3]);
  buf B_DRPADDR4 (DRPADDR_IN[4], DRPADDR[4]);
  buf B_DRPADDR5 (DRPADDR_IN[5], DRPADDR[5]);
  buf B_DRPADDR6 (DRPADDR_IN[6], DRPADDR[6]);
  buf B_DRPADDR7 (DRPADDR_IN[7], DRPADDR[7]);
  buf B_DRPADDR8 (DRPADDR_IN[8], DRPADDR[8]);
  buf B_DRPADDR9 (DRPADDR_IN[9], DRPADDR[9]);
  buf B_DRPCLK (DRPCLK_IN, DRPCLK);
  buf B_DRPDI0 (DRPDI_IN[0], DRPDI[0]);
  buf B_DRPDI1 (DRPDI_IN[1], DRPDI[1]);
  buf B_DRPDI10 (DRPDI_IN[10], DRPDI[10]);
  buf B_DRPDI11 (DRPDI_IN[11], DRPDI[11]);
  buf B_DRPDI12 (DRPDI_IN[12], DRPDI[12]);
  buf B_DRPDI13 (DRPDI_IN[13], DRPDI[13]);
  buf B_DRPDI14 (DRPDI_IN[14], DRPDI[14]);
  buf B_DRPDI15 (DRPDI_IN[15], DRPDI[15]);
  buf B_DRPDI2 (DRPDI_IN[2], DRPDI[2]);
  buf B_DRPDI3 (DRPDI_IN[3], DRPDI[3]);
  buf B_DRPDI4 (DRPDI_IN[4], DRPDI[4]);
  buf B_DRPDI5 (DRPDI_IN[5], DRPDI[5]);
  buf B_DRPDI6 (DRPDI_IN[6], DRPDI[6]);
  buf B_DRPDI7 (DRPDI_IN[7], DRPDI[7]);
  buf B_DRPDI8 (DRPDI_IN[8], DRPDI[8]);
  buf B_DRPDI9 (DRPDI_IN[9], DRPDI[9]);
  buf B_DRPEN (DRPEN_IN, DRPEN);
  buf B_DRPWE (DRPWE_IN, DRPWE);
  buf B_MAXISCQTREADY0 (MAXISCQTREADY_IN[0], MAXISCQTREADY[0]);
  buf B_MAXISCQTREADY1 (MAXISCQTREADY_IN[1], MAXISCQTREADY[1]);
  buf B_MAXISCQTREADY10 (MAXISCQTREADY_IN[10], MAXISCQTREADY[10]);
  buf B_MAXISCQTREADY11 (MAXISCQTREADY_IN[11], MAXISCQTREADY[11]);
  buf B_MAXISCQTREADY12 (MAXISCQTREADY_IN[12], MAXISCQTREADY[12]);
  buf B_MAXISCQTREADY13 (MAXISCQTREADY_IN[13], MAXISCQTREADY[13]);
  buf B_MAXISCQTREADY14 (MAXISCQTREADY_IN[14], MAXISCQTREADY[14]);
  buf B_MAXISCQTREADY15 (MAXISCQTREADY_IN[15], MAXISCQTREADY[15]);
  buf B_MAXISCQTREADY16 (MAXISCQTREADY_IN[16], MAXISCQTREADY[16]);
  buf B_MAXISCQTREADY17 (MAXISCQTREADY_IN[17], MAXISCQTREADY[17]);
  buf B_MAXISCQTREADY18 (MAXISCQTREADY_IN[18], MAXISCQTREADY[18]);
  buf B_MAXISCQTREADY19 (MAXISCQTREADY_IN[19], MAXISCQTREADY[19]);
  buf B_MAXISCQTREADY2 (MAXISCQTREADY_IN[2], MAXISCQTREADY[2]);
  buf B_MAXISCQTREADY20 (MAXISCQTREADY_IN[20], MAXISCQTREADY[20]);
  buf B_MAXISCQTREADY21 (MAXISCQTREADY_IN[21], MAXISCQTREADY[21]);
  buf B_MAXISCQTREADY3 (MAXISCQTREADY_IN[3], MAXISCQTREADY[3]);
  buf B_MAXISCQTREADY4 (MAXISCQTREADY_IN[4], MAXISCQTREADY[4]);
  buf B_MAXISCQTREADY5 (MAXISCQTREADY_IN[5], MAXISCQTREADY[5]);
  buf B_MAXISCQTREADY6 (MAXISCQTREADY_IN[6], MAXISCQTREADY[6]);
  buf B_MAXISCQTREADY7 (MAXISCQTREADY_IN[7], MAXISCQTREADY[7]);
  buf B_MAXISCQTREADY8 (MAXISCQTREADY_IN[8], MAXISCQTREADY[8]);
  buf B_MAXISCQTREADY9 (MAXISCQTREADY_IN[9], MAXISCQTREADY[9]);
  buf B_MAXISRCTREADY0 (MAXISRCTREADY_IN[0], MAXISRCTREADY[0]);
  buf B_MAXISRCTREADY1 (MAXISRCTREADY_IN[1], MAXISRCTREADY[1]);
  buf B_MAXISRCTREADY10 (MAXISRCTREADY_IN[10], MAXISRCTREADY[10]);
  buf B_MAXISRCTREADY11 (MAXISRCTREADY_IN[11], MAXISRCTREADY[11]);
  buf B_MAXISRCTREADY12 (MAXISRCTREADY_IN[12], MAXISRCTREADY[12]);
  buf B_MAXISRCTREADY13 (MAXISRCTREADY_IN[13], MAXISRCTREADY[13]);
  buf B_MAXISRCTREADY14 (MAXISRCTREADY_IN[14], MAXISRCTREADY[14]);
  buf B_MAXISRCTREADY15 (MAXISRCTREADY_IN[15], MAXISRCTREADY[15]);
  buf B_MAXISRCTREADY16 (MAXISRCTREADY_IN[16], MAXISRCTREADY[16]);
  buf B_MAXISRCTREADY17 (MAXISRCTREADY_IN[17], MAXISRCTREADY[17]);
  buf B_MAXISRCTREADY18 (MAXISRCTREADY_IN[18], MAXISRCTREADY[18]);
  buf B_MAXISRCTREADY19 (MAXISRCTREADY_IN[19], MAXISRCTREADY[19]);
  buf B_MAXISRCTREADY2 (MAXISRCTREADY_IN[2], MAXISRCTREADY[2]);
  buf B_MAXISRCTREADY20 (MAXISRCTREADY_IN[20], MAXISRCTREADY[20]);
  buf B_MAXISRCTREADY21 (MAXISRCTREADY_IN[21], MAXISRCTREADY[21]);
  buf B_MAXISRCTREADY3 (MAXISRCTREADY_IN[3], MAXISRCTREADY[3]);
  buf B_MAXISRCTREADY4 (MAXISRCTREADY_IN[4], MAXISRCTREADY[4]);
  buf B_MAXISRCTREADY5 (MAXISRCTREADY_IN[5], MAXISRCTREADY[5]);
  buf B_MAXISRCTREADY6 (MAXISRCTREADY_IN[6], MAXISRCTREADY[6]);
  buf B_MAXISRCTREADY7 (MAXISRCTREADY_IN[7], MAXISRCTREADY[7]);
  buf B_MAXISRCTREADY8 (MAXISRCTREADY_IN[8], MAXISRCTREADY[8]);
  buf B_MAXISRCTREADY9 (MAXISRCTREADY_IN[9], MAXISRCTREADY[9]);
  buf B_MGMTRESETN (MGMTRESETN_IN, MGMTRESETN);
  buf B_MGMTSTICKYRESETN (MGMTSTICKYRESETN_IN, MGMTSTICKYRESETN);
  buf B_MICOMPLETIONRAMREADDATA0 (MICOMPLETIONRAMREADDATA_IN[0], MICOMPLETIONRAMREADDATA[0]);
  buf B_MICOMPLETIONRAMREADDATA1 (MICOMPLETIONRAMREADDATA_IN[1], MICOMPLETIONRAMREADDATA[1]);
  buf B_MICOMPLETIONRAMREADDATA10 (MICOMPLETIONRAMREADDATA_IN[10], MICOMPLETIONRAMREADDATA[10]);
  buf B_MICOMPLETIONRAMREADDATA100 (MICOMPLETIONRAMREADDATA_IN[100], MICOMPLETIONRAMREADDATA[100]);
  buf B_MICOMPLETIONRAMREADDATA101 (MICOMPLETIONRAMREADDATA_IN[101], MICOMPLETIONRAMREADDATA[101]);
  buf B_MICOMPLETIONRAMREADDATA102 (MICOMPLETIONRAMREADDATA_IN[102], MICOMPLETIONRAMREADDATA[102]);
  buf B_MICOMPLETIONRAMREADDATA103 (MICOMPLETIONRAMREADDATA_IN[103], MICOMPLETIONRAMREADDATA[103]);
  buf B_MICOMPLETIONRAMREADDATA104 (MICOMPLETIONRAMREADDATA_IN[104], MICOMPLETIONRAMREADDATA[104]);
  buf B_MICOMPLETIONRAMREADDATA105 (MICOMPLETIONRAMREADDATA_IN[105], MICOMPLETIONRAMREADDATA[105]);
  buf B_MICOMPLETIONRAMREADDATA106 (MICOMPLETIONRAMREADDATA_IN[106], MICOMPLETIONRAMREADDATA[106]);
  buf B_MICOMPLETIONRAMREADDATA107 (MICOMPLETIONRAMREADDATA_IN[107], MICOMPLETIONRAMREADDATA[107]);
  buf B_MICOMPLETIONRAMREADDATA108 (MICOMPLETIONRAMREADDATA_IN[108], MICOMPLETIONRAMREADDATA[108]);
  buf B_MICOMPLETIONRAMREADDATA109 (MICOMPLETIONRAMREADDATA_IN[109], MICOMPLETIONRAMREADDATA[109]);
  buf B_MICOMPLETIONRAMREADDATA11 (MICOMPLETIONRAMREADDATA_IN[11], MICOMPLETIONRAMREADDATA[11]);
  buf B_MICOMPLETIONRAMREADDATA110 (MICOMPLETIONRAMREADDATA_IN[110], MICOMPLETIONRAMREADDATA[110]);
  buf B_MICOMPLETIONRAMREADDATA111 (MICOMPLETIONRAMREADDATA_IN[111], MICOMPLETIONRAMREADDATA[111]);
  buf B_MICOMPLETIONRAMREADDATA112 (MICOMPLETIONRAMREADDATA_IN[112], MICOMPLETIONRAMREADDATA[112]);
  buf B_MICOMPLETIONRAMREADDATA113 (MICOMPLETIONRAMREADDATA_IN[113], MICOMPLETIONRAMREADDATA[113]);
  buf B_MICOMPLETIONRAMREADDATA114 (MICOMPLETIONRAMREADDATA_IN[114], MICOMPLETIONRAMREADDATA[114]);
  buf B_MICOMPLETIONRAMREADDATA115 (MICOMPLETIONRAMREADDATA_IN[115], MICOMPLETIONRAMREADDATA[115]);
  buf B_MICOMPLETIONRAMREADDATA116 (MICOMPLETIONRAMREADDATA_IN[116], MICOMPLETIONRAMREADDATA[116]);
  buf B_MICOMPLETIONRAMREADDATA117 (MICOMPLETIONRAMREADDATA_IN[117], MICOMPLETIONRAMREADDATA[117]);
  buf B_MICOMPLETIONRAMREADDATA118 (MICOMPLETIONRAMREADDATA_IN[118], MICOMPLETIONRAMREADDATA[118]);
  buf B_MICOMPLETIONRAMREADDATA119 (MICOMPLETIONRAMREADDATA_IN[119], MICOMPLETIONRAMREADDATA[119]);
  buf B_MICOMPLETIONRAMREADDATA12 (MICOMPLETIONRAMREADDATA_IN[12], MICOMPLETIONRAMREADDATA[12]);
  buf B_MICOMPLETIONRAMREADDATA120 (MICOMPLETIONRAMREADDATA_IN[120], MICOMPLETIONRAMREADDATA[120]);
  buf B_MICOMPLETIONRAMREADDATA121 (MICOMPLETIONRAMREADDATA_IN[121], MICOMPLETIONRAMREADDATA[121]);
  buf B_MICOMPLETIONRAMREADDATA122 (MICOMPLETIONRAMREADDATA_IN[122], MICOMPLETIONRAMREADDATA[122]);
  buf B_MICOMPLETIONRAMREADDATA123 (MICOMPLETIONRAMREADDATA_IN[123], MICOMPLETIONRAMREADDATA[123]);
  buf B_MICOMPLETIONRAMREADDATA124 (MICOMPLETIONRAMREADDATA_IN[124], MICOMPLETIONRAMREADDATA[124]);
  buf B_MICOMPLETIONRAMREADDATA125 (MICOMPLETIONRAMREADDATA_IN[125], MICOMPLETIONRAMREADDATA[125]);
  buf B_MICOMPLETIONRAMREADDATA126 (MICOMPLETIONRAMREADDATA_IN[126], MICOMPLETIONRAMREADDATA[126]);
  buf B_MICOMPLETIONRAMREADDATA127 (MICOMPLETIONRAMREADDATA_IN[127], MICOMPLETIONRAMREADDATA[127]);
  buf B_MICOMPLETIONRAMREADDATA128 (MICOMPLETIONRAMREADDATA_IN[128], MICOMPLETIONRAMREADDATA[128]);
  buf B_MICOMPLETIONRAMREADDATA129 (MICOMPLETIONRAMREADDATA_IN[129], MICOMPLETIONRAMREADDATA[129]);
  buf B_MICOMPLETIONRAMREADDATA13 (MICOMPLETIONRAMREADDATA_IN[13], MICOMPLETIONRAMREADDATA[13]);
  buf B_MICOMPLETIONRAMREADDATA130 (MICOMPLETIONRAMREADDATA_IN[130], MICOMPLETIONRAMREADDATA[130]);
  buf B_MICOMPLETIONRAMREADDATA131 (MICOMPLETIONRAMREADDATA_IN[131], MICOMPLETIONRAMREADDATA[131]);
  buf B_MICOMPLETIONRAMREADDATA132 (MICOMPLETIONRAMREADDATA_IN[132], MICOMPLETIONRAMREADDATA[132]);
  buf B_MICOMPLETIONRAMREADDATA133 (MICOMPLETIONRAMREADDATA_IN[133], MICOMPLETIONRAMREADDATA[133]);
  buf B_MICOMPLETIONRAMREADDATA134 (MICOMPLETIONRAMREADDATA_IN[134], MICOMPLETIONRAMREADDATA[134]);
  buf B_MICOMPLETIONRAMREADDATA135 (MICOMPLETIONRAMREADDATA_IN[135], MICOMPLETIONRAMREADDATA[135]);
  buf B_MICOMPLETIONRAMREADDATA136 (MICOMPLETIONRAMREADDATA_IN[136], MICOMPLETIONRAMREADDATA[136]);
  buf B_MICOMPLETIONRAMREADDATA137 (MICOMPLETIONRAMREADDATA_IN[137], MICOMPLETIONRAMREADDATA[137]);
  buf B_MICOMPLETIONRAMREADDATA138 (MICOMPLETIONRAMREADDATA_IN[138], MICOMPLETIONRAMREADDATA[138]);
  buf B_MICOMPLETIONRAMREADDATA139 (MICOMPLETIONRAMREADDATA_IN[139], MICOMPLETIONRAMREADDATA[139]);
  buf B_MICOMPLETIONRAMREADDATA14 (MICOMPLETIONRAMREADDATA_IN[14], MICOMPLETIONRAMREADDATA[14]);
  buf B_MICOMPLETIONRAMREADDATA140 (MICOMPLETIONRAMREADDATA_IN[140], MICOMPLETIONRAMREADDATA[140]);
  buf B_MICOMPLETIONRAMREADDATA141 (MICOMPLETIONRAMREADDATA_IN[141], MICOMPLETIONRAMREADDATA[141]);
  buf B_MICOMPLETIONRAMREADDATA142 (MICOMPLETIONRAMREADDATA_IN[142], MICOMPLETIONRAMREADDATA[142]);
  buf B_MICOMPLETIONRAMREADDATA143 (MICOMPLETIONRAMREADDATA_IN[143], MICOMPLETIONRAMREADDATA[143]);
  buf B_MICOMPLETIONRAMREADDATA15 (MICOMPLETIONRAMREADDATA_IN[15], MICOMPLETIONRAMREADDATA[15]);
  buf B_MICOMPLETIONRAMREADDATA16 (MICOMPLETIONRAMREADDATA_IN[16], MICOMPLETIONRAMREADDATA[16]);
  buf B_MICOMPLETIONRAMREADDATA17 (MICOMPLETIONRAMREADDATA_IN[17], MICOMPLETIONRAMREADDATA[17]);
  buf B_MICOMPLETIONRAMREADDATA18 (MICOMPLETIONRAMREADDATA_IN[18], MICOMPLETIONRAMREADDATA[18]);
  buf B_MICOMPLETIONRAMREADDATA19 (MICOMPLETIONRAMREADDATA_IN[19], MICOMPLETIONRAMREADDATA[19]);
  buf B_MICOMPLETIONRAMREADDATA2 (MICOMPLETIONRAMREADDATA_IN[2], MICOMPLETIONRAMREADDATA[2]);
  buf B_MICOMPLETIONRAMREADDATA20 (MICOMPLETIONRAMREADDATA_IN[20], MICOMPLETIONRAMREADDATA[20]);
  buf B_MICOMPLETIONRAMREADDATA21 (MICOMPLETIONRAMREADDATA_IN[21], MICOMPLETIONRAMREADDATA[21]);
  buf B_MICOMPLETIONRAMREADDATA22 (MICOMPLETIONRAMREADDATA_IN[22], MICOMPLETIONRAMREADDATA[22]);
  buf B_MICOMPLETIONRAMREADDATA23 (MICOMPLETIONRAMREADDATA_IN[23], MICOMPLETIONRAMREADDATA[23]);
  buf B_MICOMPLETIONRAMREADDATA24 (MICOMPLETIONRAMREADDATA_IN[24], MICOMPLETIONRAMREADDATA[24]);
  buf B_MICOMPLETIONRAMREADDATA25 (MICOMPLETIONRAMREADDATA_IN[25], MICOMPLETIONRAMREADDATA[25]);
  buf B_MICOMPLETIONRAMREADDATA26 (MICOMPLETIONRAMREADDATA_IN[26], MICOMPLETIONRAMREADDATA[26]);
  buf B_MICOMPLETIONRAMREADDATA27 (MICOMPLETIONRAMREADDATA_IN[27], MICOMPLETIONRAMREADDATA[27]);
  buf B_MICOMPLETIONRAMREADDATA28 (MICOMPLETIONRAMREADDATA_IN[28], MICOMPLETIONRAMREADDATA[28]);
  buf B_MICOMPLETIONRAMREADDATA29 (MICOMPLETIONRAMREADDATA_IN[29], MICOMPLETIONRAMREADDATA[29]);
  buf B_MICOMPLETIONRAMREADDATA3 (MICOMPLETIONRAMREADDATA_IN[3], MICOMPLETIONRAMREADDATA[3]);
  buf B_MICOMPLETIONRAMREADDATA30 (MICOMPLETIONRAMREADDATA_IN[30], MICOMPLETIONRAMREADDATA[30]);
  buf B_MICOMPLETIONRAMREADDATA31 (MICOMPLETIONRAMREADDATA_IN[31], MICOMPLETIONRAMREADDATA[31]);
  buf B_MICOMPLETIONRAMREADDATA32 (MICOMPLETIONRAMREADDATA_IN[32], MICOMPLETIONRAMREADDATA[32]);
  buf B_MICOMPLETIONRAMREADDATA33 (MICOMPLETIONRAMREADDATA_IN[33], MICOMPLETIONRAMREADDATA[33]);
  buf B_MICOMPLETIONRAMREADDATA34 (MICOMPLETIONRAMREADDATA_IN[34], MICOMPLETIONRAMREADDATA[34]);
  buf B_MICOMPLETIONRAMREADDATA35 (MICOMPLETIONRAMREADDATA_IN[35], MICOMPLETIONRAMREADDATA[35]);
  buf B_MICOMPLETIONRAMREADDATA36 (MICOMPLETIONRAMREADDATA_IN[36], MICOMPLETIONRAMREADDATA[36]);
  buf B_MICOMPLETIONRAMREADDATA37 (MICOMPLETIONRAMREADDATA_IN[37], MICOMPLETIONRAMREADDATA[37]);
  buf B_MICOMPLETIONRAMREADDATA38 (MICOMPLETIONRAMREADDATA_IN[38], MICOMPLETIONRAMREADDATA[38]);
  buf B_MICOMPLETIONRAMREADDATA39 (MICOMPLETIONRAMREADDATA_IN[39], MICOMPLETIONRAMREADDATA[39]);
  buf B_MICOMPLETIONRAMREADDATA4 (MICOMPLETIONRAMREADDATA_IN[4], MICOMPLETIONRAMREADDATA[4]);
  buf B_MICOMPLETIONRAMREADDATA40 (MICOMPLETIONRAMREADDATA_IN[40], MICOMPLETIONRAMREADDATA[40]);
  buf B_MICOMPLETIONRAMREADDATA41 (MICOMPLETIONRAMREADDATA_IN[41], MICOMPLETIONRAMREADDATA[41]);
  buf B_MICOMPLETIONRAMREADDATA42 (MICOMPLETIONRAMREADDATA_IN[42], MICOMPLETIONRAMREADDATA[42]);
  buf B_MICOMPLETIONRAMREADDATA43 (MICOMPLETIONRAMREADDATA_IN[43], MICOMPLETIONRAMREADDATA[43]);
  buf B_MICOMPLETIONRAMREADDATA44 (MICOMPLETIONRAMREADDATA_IN[44], MICOMPLETIONRAMREADDATA[44]);
  buf B_MICOMPLETIONRAMREADDATA45 (MICOMPLETIONRAMREADDATA_IN[45], MICOMPLETIONRAMREADDATA[45]);
  buf B_MICOMPLETIONRAMREADDATA46 (MICOMPLETIONRAMREADDATA_IN[46], MICOMPLETIONRAMREADDATA[46]);
  buf B_MICOMPLETIONRAMREADDATA47 (MICOMPLETIONRAMREADDATA_IN[47], MICOMPLETIONRAMREADDATA[47]);
  buf B_MICOMPLETIONRAMREADDATA48 (MICOMPLETIONRAMREADDATA_IN[48], MICOMPLETIONRAMREADDATA[48]);
  buf B_MICOMPLETIONRAMREADDATA49 (MICOMPLETIONRAMREADDATA_IN[49], MICOMPLETIONRAMREADDATA[49]);
  buf B_MICOMPLETIONRAMREADDATA5 (MICOMPLETIONRAMREADDATA_IN[5], MICOMPLETIONRAMREADDATA[5]);
  buf B_MICOMPLETIONRAMREADDATA50 (MICOMPLETIONRAMREADDATA_IN[50], MICOMPLETIONRAMREADDATA[50]);
  buf B_MICOMPLETIONRAMREADDATA51 (MICOMPLETIONRAMREADDATA_IN[51], MICOMPLETIONRAMREADDATA[51]);
  buf B_MICOMPLETIONRAMREADDATA52 (MICOMPLETIONRAMREADDATA_IN[52], MICOMPLETIONRAMREADDATA[52]);
  buf B_MICOMPLETIONRAMREADDATA53 (MICOMPLETIONRAMREADDATA_IN[53], MICOMPLETIONRAMREADDATA[53]);
  buf B_MICOMPLETIONRAMREADDATA54 (MICOMPLETIONRAMREADDATA_IN[54], MICOMPLETIONRAMREADDATA[54]);
  buf B_MICOMPLETIONRAMREADDATA55 (MICOMPLETIONRAMREADDATA_IN[55], MICOMPLETIONRAMREADDATA[55]);
  buf B_MICOMPLETIONRAMREADDATA56 (MICOMPLETIONRAMREADDATA_IN[56], MICOMPLETIONRAMREADDATA[56]);
  buf B_MICOMPLETIONRAMREADDATA57 (MICOMPLETIONRAMREADDATA_IN[57], MICOMPLETIONRAMREADDATA[57]);
  buf B_MICOMPLETIONRAMREADDATA58 (MICOMPLETIONRAMREADDATA_IN[58], MICOMPLETIONRAMREADDATA[58]);
  buf B_MICOMPLETIONRAMREADDATA59 (MICOMPLETIONRAMREADDATA_IN[59], MICOMPLETIONRAMREADDATA[59]);
  buf B_MICOMPLETIONRAMREADDATA6 (MICOMPLETIONRAMREADDATA_IN[6], MICOMPLETIONRAMREADDATA[6]);
  buf B_MICOMPLETIONRAMREADDATA60 (MICOMPLETIONRAMREADDATA_IN[60], MICOMPLETIONRAMREADDATA[60]);
  buf B_MICOMPLETIONRAMREADDATA61 (MICOMPLETIONRAMREADDATA_IN[61], MICOMPLETIONRAMREADDATA[61]);
  buf B_MICOMPLETIONRAMREADDATA62 (MICOMPLETIONRAMREADDATA_IN[62], MICOMPLETIONRAMREADDATA[62]);
  buf B_MICOMPLETIONRAMREADDATA63 (MICOMPLETIONRAMREADDATA_IN[63], MICOMPLETIONRAMREADDATA[63]);
  buf B_MICOMPLETIONRAMREADDATA64 (MICOMPLETIONRAMREADDATA_IN[64], MICOMPLETIONRAMREADDATA[64]);
  buf B_MICOMPLETIONRAMREADDATA65 (MICOMPLETIONRAMREADDATA_IN[65], MICOMPLETIONRAMREADDATA[65]);
  buf B_MICOMPLETIONRAMREADDATA66 (MICOMPLETIONRAMREADDATA_IN[66], MICOMPLETIONRAMREADDATA[66]);
  buf B_MICOMPLETIONRAMREADDATA67 (MICOMPLETIONRAMREADDATA_IN[67], MICOMPLETIONRAMREADDATA[67]);
  buf B_MICOMPLETIONRAMREADDATA68 (MICOMPLETIONRAMREADDATA_IN[68], MICOMPLETIONRAMREADDATA[68]);
  buf B_MICOMPLETIONRAMREADDATA69 (MICOMPLETIONRAMREADDATA_IN[69], MICOMPLETIONRAMREADDATA[69]);
  buf B_MICOMPLETIONRAMREADDATA7 (MICOMPLETIONRAMREADDATA_IN[7], MICOMPLETIONRAMREADDATA[7]);
  buf B_MICOMPLETIONRAMREADDATA70 (MICOMPLETIONRAMREADDATA_IN[70], MICOMPLETIONRAMREADDATA[70]);
  buf B_MICOMPLETIONRAMREADDATA71 (MICOMPLETIONRAMREADDATA_IN[71], MICOMPLETIONRAMREADDATA[71]);
  buf B_MICOMPLETIONRAMREADDATA72 (MICOMPLETIONRAMREADDATA_IN[72], MICOMPLETIONRAMREADDATA[72]);
  buf B_MICOMPLETIONRAMREADDATA73 (MICOMPLETIONRAMREADDATA_IN[73], MICOMPLETIONRAMREADDATA[73]);
  buf B_MICOMPLETIONRAMREADDATA74 (MICOMPLETIONRAMREADDATA_IN[74], MICOMPLETIONRAMREADDATA[74]);
  buf B_MICOMPLETIONRAMREADDATA75 (MICOMPLETIONRAMREADDATA_IN[75], MICOMPLETIONRAMREADDATA[75]);
  buf B_MICOMPLETIONRAMREADDATA76 (MICOMPLETIONRAMREADDATA_IN[76], MICOMPLETIONRAMREADDATA[76]);
  buf B_MICOMPLETIONRAMREADDATA77 (MICOMPLETIONRAMREADDATA_IN[77], MICOMPLETIONRAMREADDATA[77]);
  buf B_MICOMPLETIONRAMREADDATA78 (MICOMPLETIONRAMREADDATA_IN[78], MICOMPLETIONRAMREADDATA[78]);
  buf B_MICOMPLETIONRAMREADDATA79 (MICOMPLETIONRAMREADDATA_IN[79], MICOMPLETIONRAMREADDATA[79]);
  buf B_MICOMPLETIONRAMREADDATA8 (MICOMPLETIONRAMREADDATA_IN[8], MICOMPLETIONRAMREADDATA[8]);
  buf B_MICOMPLETIONRAMREADDATA80 (MICOMPLETIONRAMREADDATA_IN[80], MICOMPLETIONRAMREADDATA[80]);
  buf B_MICOMPLETIONRAMREADDATA81 (MICOMPLETIONRAMREADDATA_IN[81], MICOMPLETIONRAMREADDATA[81]);
  buf B_MICOMPLETIONRAMREADDATA82 (MICOMPLETIONRAMREADDATA_IN[82], MICOMPLETIONRAMREADDATA[82]);
  buf B_MICOMPLETIONRAMREADDATA83 (MICOMPLETIONRAMREADDATA_IN[83], MICOMPLETIONRAMREADDATA[83]);
  buf B_MICOMPLETIONRAMREADDATA84 (MICOMPLETIONRAMREADDATA_IN[84], MICOMPLETIONRAMREADDATA[84]);
  buf B_MICOMPLETIONRAMREADDATA85 (MICOMPLETIONRAMREADDATA_IN[85], MICOMPLETIONRAMREADDATA[85]);
  buf B_MICOMPLETIONRAMREADDATA86 (MICOMPLETIONRAMREADDATA_IN[86], MICOMPLETIONRAMREADDATA[86]);
  buf B_MICOMPLETIONRAMREADDATA87 (MICOMPLETIONRAMREADDATA_IN[87], MICOMPLETIONRAMREADDATA[87]);
  buf B_MICOMPLETIONRAMREADDATA88 (MICOMPLETIONRAMREADDATA_IN[88], MICOMPLETIONRAMREADDATA[88]);
  buf B_MICOMPLETIONRAMREADDATA89 (MICOMPLETIONRAMREADDATA_IN[89], MICOMPLETIONRAMREADDATA[89]);
  buf B_MICOMPLETIONRAMREADDATA9 (MICOMPLETIONRAMREADDATA_IN[9], MICOMPLETIONRAMREADDATA[9]);
  buf B_MICOMPLETIONRAMREADDATA90 (MICOMPLETIONRAMREADDATA_IN[90], MICOMPLETIONRAMREADDATA[90]);
  buf B_MICOMPLETIONRAMREADDATA91 (MICOMPLETIONRAMREADDATA_IN[91], MICOMPLETIONRAMREADDATA[91]);
  buf B_MICOMPLETIONRAMREADDATA92 (MICOMPLETIONRAMREADDATA_IN[92], MICOMPLETIONRAMREADDATA[92]);
  buf B_MICOMPLETIONRAMREADDATA93 (MICOMPLETIONRAMREADDATA_IN[93], MICOMPLETIONRAMREADDATA[93]);
  buf B_MICOMPLETIONRAMREADDATA94 (MICOMPLETIONRAMREADDATA_IN[94], MICOMPLETIONRAMREADDATA[94]);
  buf B_MICOMPLETIONRAMREADDATA95 (MICOMPLETIONRAMREADDATA_IN[95], MICOMPLETIONRAMREADDATA[95]);
  buf B_MICOMPLETIONRAMREADDATA96 (MICOMPLETIONRAMREADDATA_IN[96], MICOMPLETIONRAMREADDATA[96]);
  buf B_MICOMPLETIONRAMREADDATA97 (MICOMPLETIONRAMREADDATA_IN[97], MICOMPLETIONRAMREADDATA[97]);
  buf B_MICOMPLETIONRAMREADDATA98 (MICOMPLETIONRAMREADDATA_IN[98], MICOMPLETIONRAMREADDATA[98]);
  buf B_MICOMPLETIONRAMREADDATA99 (MICOMPLETIONRAMREADDATA_IN[99], MICOMPLETIONRAMREADDATA[99]);
  buf B_MIREPLAYRAMREADDATA0 (MIREPLAYRAMREADDATA_IN[0], MIREPLAYRAMREADDATA[0]);
  buf B_MIREPLAYRAMREADDATA1 (MIREPLAYRAMREADDATA_IN[1], MIREPLAYRAMREADDATA[1]);
  buf B_MIREPLAYRAMREADDATA10 (MIREPLAYRAMREADDATA_IN[10], MIREPLAYRAMREADDATA[10]);
  buf B_MIREPLAYRAMREADDATA100 (MIREPLAYRAMREADDATA_IN[100], MIREPLAYRAMREADDATA[100]);
  buf B_MIREPLAYRAMREADDATA101 (MIREPLAYRAMREADDATA_IN[101], MIREPLAYRAMREADDATA[101]);
  buf B_MIREPLAYRAMREADDATA102 (MIREPLAYRAMREADDATA_IN[102], MIREPLAYRAMREADDATA[102]);
  buf B_MIREPLAYRAMREADDATA103 (MIREPLAYRAMREADDATA_IN[103], MIREPLAYRAMREADDATA[103]);
  buf B_MIREPLAYRAMREADDATA104 (MIREPLAYRAMREADDATA_IN[104], MIREPLAYRAMREADDATA[104]);
  buf B_MIREPLAYRAMREADDATA105 (MIREPLAYRAMREADDATA_IN[105], MIREPLAYRAMREADDATA[105]);
  buf B_MIREPLAYRAMREADDATA106 (MIREPLAYRAMREADDATA_IN[106], MIREPLAYRAMREADDATA[106]);
  buf B_MIREPLAYRAMREADDATA107 (MIREPLAYRAMREADDATA_IN[107], MIREPLAYRAMREADDATA[107]);
  buf B_MIREPLAYRAMREADDATA108 (MIREPLAYRAMREADDATA_IN[108], MIREPLAYRAMREADDATA[108]);
  buf B_MIREPLAYRAMREADDATA109 (MIREPLAYRAMREADDATA_IN[109], MIREPLAYRAMREADDATA[109]);
  buf B_MIREPLAYRAMREADDATA11 (MIREPLAYRAMREADDATA_IN[11], MIREPLAYRAMREADDATA[11]);
  buf B_MIREPLAYRAMREADDATA110 (MIREPLAYRAMREADDATA_IN[110], MIREPLAYRAMREADDATA[110]);
  buf B_MIREPLAYRAMREADDATA111 (MIREPLAYRAMREADDATA_IN[111], MIREPLAYRAMREADDATA[111]);
  buf B_MIREPLAYRAMREADDATA112 (MIREPLAYRAMREADDATA_IN[112], MIREPLAYRAMREADDATA[112]);
  buf B_MIREPLAYRAMREADDATA113 (MIREPLAYRAMREADDATA_IN[113], MIREPLAYRAMREADDATA[113]);
  buf B_MIREPLAYRAMREADDATA114 (MIREPLAYRAMREADDATA_IN[114], MIREPLAYRAMREADDATA[114]);
  buf B_MIREPLAYRAMREADDATA115 (MIREPLAYRAMREADDATA_IN[115], MIREPLAYRAMREADDATA[115]);
  buf B_MIREPLAYRAMREADDATA116 (MIREPLAYRAMREADDATA_IN[116], MIREPLAYRAMREADDATA[116]);
  buf B_MIREPLAYRAMREADDATA117 (MIREPLAYRAMREADDATA_IN[117], MIREPLAYRAMREADDATA[117]);
  buf B_MIREPLAYRAMREADDATA118 (MIREPLAYRAMREADDATA_IN[118], MIREPLAYRAMREADDATA[118]);
  buf B_MIREPLAYRAMREADDATA119 (MIREPLAYRAMREADDATA_IN[119], MIREPLAYRAMREADDATA[119]);
  buf B_MIREPLAYRAMREADDATA12 (MIREPLAYRAMREADDATA_IN[12], MIREPLAYRAMREADDATA[12]);
  buf B_MIREPLAYRAMREADDATA120 (MIREPLAYRAMREADDATA_IN[120], MIREPLAYRAMREADDATA[120]);
  buf B_MIREPLAYRAMREADDATA121 (MIREPLAYRAMREADDATA_IN[121], MIREPLAYRAMREADDATA[121]);
  buf B_MIREPLAYRAMREADDATA122 (MIREPLAYRAMREADDATA_IN[122], MIREPLAYRAMREADDATA[122]);
  buf B_MIREPLAYRAMREADDATA123 (MIREPLAYRAMREADDATA_IN[123], MIREPLAYRAMREADDATA[123]);
  buf B_MIREPLAYRAMREADDATA124 (MIREPLAYRAMREADDATA_IN[124], MIREPLAYRAMREADDATA[124]);
  buf B_MIREPLAYRAMREADDATA125 (MIREPLAYRAMREADDATA_IN[125], MIREPLAYRAMREADDATA[125]);
  buf B_MIREPLAYRAMREADDATA126 (MIREPLAYRAMREADDATA_IN[126], MIREPLAYRAMREADDATA[126]);
  buf B_MIREPLAYRAMREADDATA127 (MIREPLAYRAMREADDATA_IN[127], MIREPLAYRAMREADDATA[127]);
  buf B_MIREPLAYRAMREADDATA128 (MIREPLAYRAMREADDATA_IN[128], MIREPLAYRAMREADDATA[128]);
  buf B_MIREPLAYRAMREADDATA129 (MIREPLAYRAMREADDATA_IN[129], MIREPLAYRAMREADDATA[129]);
  buf B_MIREPLAYRAMREADDATA13 (MIREPLAYRAMREADDATA_IN[13], MIREPLAYRAMREADDATA[13]);
  buf B_MIREPLAYRAMREADDATA130 (MIREPLAYRAMREADDATA_IN[130], MIREPLAYRAMREADDATA[130]);
  buf B_MIREPLAYRAMREADDATA131 (MIREPLAYRAMREADDATA_IN[131], MIREPLAYRAMREADDATA[131]);
  buf B_MIREPLAYRAMREADDATA132 (MIREPLAYRAMREADDATA_IN[132], MIREPLAYRAMREADDATA[132]);
  buf B_MIREPLAYRAMREADDATA133 (MIREPLAYRAMREADDATA_IN[133], MIREPLAYRAMREADDATA[133]);
  buf B_MIREPLAYRAMREADDATA134 (MIREPLAYRAMREADDATA_IN[134], MIREPLAYRAMREADDATA[134]);
  buf B_MIREPLAYRAMREADDATA135 (MIREPLAYRAMREADDATA_IN[135], MIREPLAYRAMREADDATA[135]);
  buf B_MIREPLAYRAMREADDATA136 (MIREPLAYRAMREADDATA_IN[136], MIREPLAYRAMREADDATA[136]);
  buf B_MIREPLAYRAMREADDATA137 (MIREPLAYRAMREADDATA_IN[137], MIREPLAYRAMREADDATA[137]);
  buf B_MIREPLAYRAMREADDATA138 (MIREPLAYRAMREADDATA_IN[138], MIREPLAYRAMREADDATA[138]);
  buf B_MIREPLAYRAMREADDATA139 (MIREPLAYRAMREADDATA_IN[139], MIREPLAYRAMREADDATA[139]);
  buf B_MIREPLAYRAMREADDATA14 (MIREPLAYRAMREADDATA_IN[14], MIREPLAYRAMREADDATA[14]);
  buf B_MIREPLAYRAMREADDATA140 (MIREPLAYRAMREADDATA_IN[140], MIREPLAYRAMREADDATA[140]);
  buf B_MIREPLAYRAMREADDATA141 (MIREPLAYRAMREADDATA_IN[141], MIREPLAYRAMREADDATA[141]);
  buf B_MIREPLAYRAMREADDATA142 (MIREPLAYRAMREADDATA_IN[142], MIREPLAYRAMREADDATA[142]);
  buf B_MIREPLAYRAMREADDATA143 (MIREPLAYRAMREADDATA_IN[143], MIREPLAYRAMREADDATA[143]);
  buf B_MIREPLAYRAMREADDATA15 (MIREPLAYRAMREADDATA_IN[15], MIREPLAYRAMREADDATA[15]);
  buf B_MIREPLAYRAMREADDATA16 (MIREPLAYRAMREADDATA_IN[16], MIREPLAYRAMREADDATA[16]);
  buf B_MIREPLAYRAMREADDATA17 (MIREPLAYRAMREADDATA_IN[17], MIREPLAYRAMREADDATA[17]);
  buf B_MIREPLAYRAMREADDATA18 (MIREPLAYRAMREADDATA_IN[18], MIREPLAYRAMREADDATA[18]);
  buf B_MIREPLAYRAMREADDATA19 (MIREPLAYRAMREADDATA_IN[19], MIREPLAYRAMREADDATA[19]);
  buf B_MIREPLAYRAMREADDATA2 (MIREPLAYRAMREADDATA_IN[2], MIREPLAYRAMREADDATA[2]);
  buf B_MIREPLAYRAMREADDATA20 (MIREPLAYRAMREADDATA_IN[20], MIREPLAYRAMREADDATA[20]);
  buf B_MIREPLAYRAMREADDATA21 (MIREPLAYRAMREADDATA_IN[21], MIREPLAYRAMREADDATA[21]);
  buf B_MIREPLAYRAMREADDATA22 (MIREPLAYRAMREADDATA_IN[22], MIREPLAYRAMREADDATA[22]);
  buf B_MIREPLAYRAMREADDATA23 (MIREPLAYRAMREADDATA_IN[23], MIREPLAYRAMREADDATA[23]);
  buf B_MIREPLAYRAMREADDATA24 (MIREPLAYRAMREADDATA_IN[24], MIREPLAYRAMREADDATA[24]);
  buf B_MIREPLAYRAMREADDATA25 (MIREPLAYRAMREADDATA_IN[25], MIREPLAYRAMREADDATA[25]);
  buf B_MIREPLAYRAMREADDATA26 (MIREPLAYRAMREADDATA_IN[26], MIREPLAYRAMREADDATA[26]);
  buf B_MIREPLAYRAMREADDATA27 (MIREPLAYRAMREADDATA_IN[27], MIREPLAYRAMREADDATA[27]);
  buf B_MIREPLAYRAMREADDATA28 (MIREPLAYRAMREADDATA_IN[28], MIREPLAYRAMREADDATA[28]);
  buf B_MIREPLAYRAMREADDATA29 (MIREPLAYRAMREADDATA_IN[29], MIREPLAYRAMREADDATA[29]);
  buf B_MIREPLAYRAMREADDATA3 (MIREPLAYRAMREADDATA_IN[3], MIREPLAYRAMREADDATA[3]);
  buf B_MIREPLAYRAMREADDATA30 (MIREPLAYRAMREADDATA_IN[30], MIREPLAYRAMREADDATA[30]);
  buf B_MIREPLAYRAMREADDATA31 (MIREPLAYRAMREADDATA_IN[31], MIREPLAYRAMREADDATA[31]);
  buf B_MIREPLAYRAMREADDATA32 (MIREPLAYRAMREADDATA_IN[32], MIREPLAYRAMREADDATA[32]);
  buf B_MIREPLAYRAMREADDATA33 (MIREPLAYRAMREADDATA_IN[33], MIREPLAYRAMREADDATA[33]);
  buf B_MIREPLAYRAMREADDATA34 (MIREPLAYRAMREADDATA_IN[34], MIREPLAYRAMREADDATA[34]);
  buf B_MIREPLAYRAMREADDATA35 (MIREPLAYRAMREADDATA_IN[35], MIREPLAYRAMREADDATA[35]);
  buf B_MIREPLAYRAMREADDATA36 (MIREPLAYRAMREADDATA_IN[36], MIREPLAYRAMREADDATA[36]);
  buf B_MIREPLAYRAMREADDATA37 (MIREPLAYRAMREADDATA_IN[37], MIREPLAYRAMREADDATA[37]);
  buf B_MIREPLAYRAMREADDATA38 (MIREPLAYRAMREADDATA_IN[38], MIREPLAYRAMREADDATA[38]);
  buf B_MIREPLAYRAMREADDATA39 (MIREPLAYRAMREADDATA_IN[39], MIREPLAYRAMREADDATA[39]);
  buf B_MIREPLAYRAMREADDATA4 (MIREPLAYRAMREADDATA_IN[4], MIREPLAYRAMREADDATA[4]);
  buf B_MIREPLAYRAMREADDATA40 (MIREPLAYRAMREADDATA_IN[40], MIREPLAYRAMREADDATA[40]);
  buf B_MIREPLAYRAMREADDATA41 (MIREPLAYRAMREADDATA_IN[41], MIREPLAYRAMREADDATA[41]);
  buf B_MIREPLAYRAMREADDATA42 (MIREPLAYRAMREADDATA_IN[42], MIREPLAYRAMREADDATA[42]);
  buf B_MIREPLAYRAMREADDATA43 (MIREPLAYRAMREADDATA_IN[43], MIREPLAYRAMREADDATA[43]);
  buf B_MIREPLAYRAMREADDATA44 (MIREPLAYRAMREADDATA_IN[44], MIREPLAYRAMREADDATA[44]);
  buf B_MIREPLAYRAMREADDATA45 (MIREPLAYRAMREADDATA_IN[45], MIREPLAYRAMREADDATA[45]);
  buf B_MIREPLAYRAMREADDATA46 (MIREPLAYRAMREADDATA_IN[46], MIREPLAYRAMREADDATA[46]);
  buf B_MIREPLAYRAMREADDATA47 (MIREPLAYRAMREADDATA_IN[47], MIREPLAYRAMREADDATA[47]);
  buf B_MIREPLAYRAMREADDATA48 (MIREPLAYRAMREADDATA_IN[48], MIREPLAYRAMREADDATA[48]);
  buf B_MIREPLAYRAMREADDATA49 (MIREPLAYRAMREADDATA_IN[49], MIREPLAYRAMREADDATA[49]);
  buf B_MIREPLAYRAMREADDATA5 (MIREPLAYRAMREADDATA_IN[5], MIREPLAYRAMREADDATA[5]);
  buf B_MIREPLAYRAMREADDATA50 (MIREPLAYRAMREADDATA_IN[50], MIREPLAYRAMREADDATA[50]);
  buf B_MIREPLAYRAMREADDATA51 (MIREPLAYRAMREADDATA_IN[51], MIREPLAYRAMREADDATA[51]);
  buf B_MIREPLAYRAMREADDATA52 (MIREPLAYRAMREADDATA_IN[52], MIREPLAYRAMREADDATA[52]);
  buf B_MIREPLAYRAMREADDATA53 (MIREPLAYRAMREADDATA_IN[53], MIREPLAYRAMREADDATA[53]);
  buf B_MIREPLAYRAMREADDATA54 (MIREPLAYRAMREADDATA_IN[54], MIREPLAYRAMREADDATA[54]);
  buf B_MIREPLAYRAMREADDATA55 (MIREPLAYRAMREADDATA_IN[55], MIREPLAYRAMREADDATA[55]);
  buf B_MIREPLAYRAMREADDATA56 (MIREPLAYRAMREADDATA_IN[56], MIREPLAYRAMREADDATA[56]);
  buf B_MIREPLAYRAMREADDATA57 (MIREPLAYRAMREADDATA_IN[57], MIREPLAYRAMREADDATA[57]);
  buf B_MIREPLAYRAMREADDATA58 (MIREPLAYRAMREADDATA_IN[58], MIREPLAYRAMREADDATA[58]);
  buf B_MIREPLAYRAMREADDATA59 (MIREPLAYRAMREADDATA_IN[59], MIREPLAYRAMREADDATA[59]);
  buf B_MIREPLAYRAMREADDATA6 (MIREPLAYRAMREADDATA_IN[6], MIREPLAYRAMREADDATA[6]);
  buf B_MIREPLAYRAMREADDATA60 (MIREPLAYRAMREADDATA_IN[60], MIREPLAYRAMREADDATA[60]);
  buf B_MIREPLAYRAMREADDATA61 (MIREPLAYRAMREADDATA_IN[61], MIREPLAYRAMREADDATA[61]);
  buf B_MIREPLAYRAMREADDATA62 (MIREPLAYRAMREADDATA_IN[62], MIREPLAYRAMREADDATA[62]);
  buf B_MIREPLAYRAMREADDATA63 (MIREPLAYRAMREADDATA_IN[63], MIREPLAYRAMREADDATA[63]);
  buf B_MIREPLAYRAMREADDATA64 (MIREPLAYRAMREADDATA_IN[64], MIREPLAYRAMREADDATA[64]);
  buf B_MIREPLAYRAMREADDATA65 (MIREPLAYRAMREADDATA_IN[65], MIREPLAYRAMREADDATA[65]);
  buf B_MIREPLAYRAMREADDATA66 (MIREPLAYRAMREADDATA_IN[66], MIREPLAYRAMREADDATA[66]);
  buf B_MIREPLAYRAMREADDATA67 (MIREPLAYRAMREADDATA_IN[67], MIREPLAYRAMREADDATA[67]);
  buf B_MIREPLAYRAMREADDATA68 (MIREPLAYRAMREADDATA_IN[68], MIREPLAYRAMREADDATA[68]);
  buf B_MIREPLAYRAMREADDATA69 (MIREPLAYRAMREADDATA_IN[69], MIREPLAYRAMREADDATA[69]);
  buf B_MIREPLAYRAMREADDATA7 (MIREPLAYRAMREADDATA_IN[7], MIREPLAYRAMREADDATA[7]);
  buf B_MIREPLAYRAMREADDATA70 (MIREPLAYRAMREADDATA_IN[70], MIREPLAYRAMREADDATA[70]);
  buf B_MIREPLAYRAMREADDATA71 (MIREPLAYRAMREADDATA_IN[71], MIREPLAYRAMREADDATA[71]);
  buf B_MIREPLAYRAMREADDATA72 (MIREPLAYRAMREADDATA_IN[72], MIREPLAYRAMREADDATA[72]);
  buf B_MIREPLAYRAMREADDATA73 (MIREPLAYRAMREADDATA_IN[73], MIREPLAYRAMREADDATA[73]);
  buf B_MIREPLAYRAMREADDATA74 (MIREPLAYRAMREADDATA_IN[74], MIREPLAYRAMREADDATA[74]);
  buf B_MIREPLAYRAMREADDATA75 (MIREPLAYRAMREADDATA_IN[75], MIREPLAYRAMREADDATA[75]);
  buf B_MIREPLAYRAMREADDATA76 (MIREPLAYRAMREADDATA_IN[76], MIREPLAYRAMREADDATA[76]);
  buf B_MIREPLAYRAMREADDATA77 (MIREPLAYRAMREADDATA_IN[77], MIREPLAYRAMREADDATA[77]);
  buf B_MIREPLAYRAMREADDATA78 (MIREPLAYRAMREADDATA_IN[78], MIREPLAYRAMREADDATA[78]);
  buf B_MIREPLAYRAMREADDATA79 (MIREPLAYRAMREADDATA_IN[79], MIREPLAYRAMREADDATA[79]);
  buf B_MIREPLAYRAMREADDATA8 (MIREPLAYRAMREADDATA_IN[8], MIREPLAYRAMREADDATA[8]);
  buf B_MIREPLAYRAMREADDATA80 (MIREPLAYRAMREADDATA_IN[80], MIREPLAYRAMREADDATA[80]);
  buf B_MIREPLAYRAMREADDATA81 (MIREPLAYRAMREADDATA_IN[81], MIREPLAYRAMREADDATA[81]);
  buf B_MIREPLAYRAMREADDATA82 (MIREPLAYRAMREADDATA_IN[82], MIREPLAYRAMREADDATA[82]);
  buf B_MIREPLAYRAMREADDATA83 (MIREPLAYRAMREADDATA_IN[83], MIREPLAYRAMREADDATA[83]);
  buf B_MIREPLAYRAMREADDATA84 (MIREPLAYRAMREADDATA_IN[84], MIREPLAYRAMREADDATA[84]);
  buf B_MIREPLAYRAMREADDATA85 (MIREPLAYRAMREADDATA_IN[85], MIREPLAYRAMREADDATA[85]);
  buf B_MIREPLAYRAMREADDATA86 (MIREPLAYRAMREADDATA_IN[86], MIREPLAYRAMREADDATA[86]);
  buf B_MIREPLAYRAMREADDATA87 (MIREPLAYRAMREADDATA_IN[87], MIREPLAYRAMREADDATA[87]);
  buf B_MIREPLAYRAMREADDATA88 (MIREPLAYRAMREADDATA_IN[88], MIREPLAYRAMREADDATA[88]);
  buf B_MIREPLAYRAMREADDATA89 (MIREPLAYRAMREADDATA_IN[89], MIREPLAYRAMREADDATA[89]);
  buf B_MIREPLAYRAMREADDATA9 (MIREPLAYRAMREADDATA_IN[9], MIREPLAYRAMREADDATA[9]);
  buf B_MIREPLAYRAMREADDATA90 (MIREPLAYRAMREADDATA_IN[90], MIREPLAYRAMREADDATA[90]);
  buf B_MIREPLAYRAMREADDATA91 (MIREPLAYRAMREADDATA_IN[91], MIREPLAYRAMREADDATA[91]);
  buf B_MIREPLAYRAMREADDATA92 (MIREPLAYRAMREADDATA_IN[92], MIREPLAYRAMREADDATA[92]);
  buf B_MIREPLAYRAMREADDATA93 (MIREPLAYRAMREADDATA_IN[93], MIREPLAYRAMREADDATA[93]);
  buf B_MIREPLAYRAMREADDATA94 (MIREPLAYRAMREADDATA_IN[94], MIREPLAYRAMREADDATA[94]);
  buf B_MIREPLAYRAMREADDATA95 (MIREPLAYRAMREADDATA_IN[95], MIREPLAYRAMREADDATA[95]);
  buf B_MIREPLAYRAMREADDATA96 (MIREPLAYRAMREADDATA_IN[96], MIREPLAYRAMREADDATA[96]);
  buf B_MIREPLAYRAMREADDATA97 (MIREPLAYRAMREADDATA_IN[97], MIREPLAYRAMREADDATA[97]);
  buf B_MIREPLAYRAMREADDATA98 (MIREPLAYRAMREADDATA_IN[98], MIREPLAYRAMREADDATA[98]);
  buf B_MIREPLAYRAMREADDATA99 (MIREPLAYRAMREADDATA_IN[99], MIREPLAYRAMREADDATA[99]);
  buf B_MIREQUESTRAMREADDATA0 (MIREQUESTRAMREADDATA_IN[0], MIREQUESTRAMREADDATA[0]);
  buf B_MIREQUESTRAMREADDATA1 (MIREQUESTRAMREADDATA_IN[1], MIREQUESTRAMREADDATA[1]);
  buf B_MIREQUESTRAMREADDATA10 (MIREQUESTRAMREADDATA_IN[10], MIREQUESTRAMREADDATA[10]);
  buf B_MIREQUESTRAMREADDATA100 (MIREQUESTRAMREADDATA_IN[100], MIREQUESTRAMREADDATA[100]);
  buf B_MIREQUESTRAMREADDATA101 (MIREQUESTRAMREADDATA_IN[101], MIREQUESTRAMREADDATA[101]);
  buf B_MIREQUESTRAMREADDATA102 (MIREQUESTRAMREADDATA_IN[102], MIREQUESTRAMREADDATA[102]);
  buf B_MIREQUESTRAMREADDATA103 (MIREQUESTRAMREADDATA_IN[103], MIREQUESTRAMREADDATA[103]);
  buf B_MIREQUESTRAMREADDATA104 (MIREQUESTRAMREADDATA_IN[104], MIREQUESTRAMREADDATA[104]);
  buf B_MIREQUESTRAMREADDATA105 (MIREQUESTRAMREADDATA_IN[105], MIREQUESTRAMREADDATA[105]);
  buf B_MIREQUESTRAMREADDATA106 (MIREQUESTRAMREADDATA_IN[106], MIREQUESTRAMREADDATA[106]);
  buf B_MIREQUESTRAMREADDATA107 (MIREQUESTRAMREADDATA_IN[107], MIREQUESTRAMREADDATA[107]);
  buf B_MIREQUESTRAMREADDATA108 (MIREQUESTRAMREADDATA_IN[108], MIREQUESTRAMREADDATA[108]);
  buf B_MIREQUESTRAMREADDATA109 (MIREQUESTRAMREADDATA_IN[109], MIREQUESTRAMREADDATA[109]);
  buf B_MIREQUESTRAMREADDATA11 (MIREQUESTRAMREADDATA_IN[11], MIREQUESTRAMREADDATA[11]);
  buf B_MIREQUESTRAMREADDATA110 (MIREQUESTRAMREADDATA_IN[110], MIREQUESTRAMREADDATA[110]);
  buf B_MIREQUESTRAMREADDATA111 (MIREQUESTRAMREADDATA_IN[111], MIREQUESTRAMREADDATA[111]);
  buf B_MIREQUESTRAMREADDATA112 (MIREQUESTRAMREADDATA_IN[112], MIREQUESTRAMREADDATA[112]);
  buf B_MIREQUESTRAMREADDATA113 (MIREQUESTRAMREADDATA_IN[113], MIREQUESTRAMREADDATA[113]);
  buf B_MIREQUESTRAMREADDATA114 (MIREQUESTRAMREADDATA_IN[114], MIREQUESTRAMREADDATA[114]);
  buf B_MIREQUESTRAMREADDATA115 (MIREQUESTRAMREADDATA_IN[115], MIREQUESTRAMREADDATA[115]);
  buf B_MIREQUESTRAMREADDATA116 (MIREQUESTRAMREADDATA_IN[116], MIREQUESTRAMREADDATA[116]);
  buf B_MIREQUESTRAMREADDATA117 (MIREQUESTRAMREADDATA_IN[117], MIREQUESTRAMREADDATA[117]);
  buf B_MIREQUESTRAMREADDATA118 (MIREQUESTRAMREADDATA_IN[118], MIREQUESTRAMREADDATA[118]);
  buf B_MIREQUESTRAMREADDATA119 (MIREQUESTRAMREADDATA_IN[119], MIREQUESTRAMREADDATA[119]);
  buf B_MIREQUESTRAMREADDATA12 (MIREQUESTRAMREADDATA_IN[12], MIREQUESTRAMREADDATA[12]);
  buf B_MIREQUESTRAMREADDATA120 (MIREQUESTRAMREADDATA_IN[120], MIREQUESTRAMREADDATA[120]);
  buf B_MIREQUESTRAMREADDATA121 (MIREQUESTRAMREADDATA_IN[121], MIREQUESTRAMREADDATA[121]);
  buf B_MIREQUESTRAMREADDATA122 (MIREQUESTRAMREADDATA_IN[122], MIREQUESTRAMREADDATA[122]);
  buf B_MIREQUESTRAMREADDATA123 (MIREQUESTRAMREADDATA_IN[123], MIREQUESTRAMREADDATA[123]);
  buf B_MIREQUESTRAMREADDATA124 (MIREQUESTRAMREADDATA_IN[124], MIREQUESTRAMREADDATA[124]);
  buf B_MIREQUESTRAMREADDATA125 (MIREQUESTRAMREADDATA_IN[125], MIREQUESTRAMREADDATA[125]);
  buf B_MIREQUESTRAMREADDATA126 (MIREQUESTRAMREADDATA_IN[126], MIREQUESTRAMREADDATA[126]);
  buf B_MIREQUESTRAMREADDATA127 (MIREQUESTRAMREADDATA_IN[127], MIREQUESTRAMREADDATA[127]);
  buf B_MIREQUESTRAMREADDATA128 (MIREQUESTRAMREADDATA_IN[128], MIREQUESTRAMREADDATA[128]);
  buf B_MIREQUESTRAMREADDATA129 (MIREQUESTRAMREADDATA_IN[129], MIREQUESTRAMREADDATA[129]);
  buf B_MIREQUESTRAMREADDATA13 (MIREQUESTRAMREADDATA_IN[13], MIREQUESTRAMREADDATA[13]);
  buf B_MIREQUESTRAMREADDATA130 (MIREQUESTRAMREADDATA_IN[130], MIREQUESTRAMREADDATA[130]);
  buf B_MIREQUESTRAMREADDATA131 (MIREQUESTRAMREADDATA_IN[131], MIREQUESTRAMREADDATA[131]);
  buf B_MIREQUESTRAMREADDATA132 (MIREQUESTRAMREADDATA_IN[132], MIREQUESTRAMREADDATA[132]);
  buf B_MIREQUESTRAMREADDATA133 (MIREQUESTRAMREADDATA_IN[133], MIREQUESTRAMREADDATA[133]);
  buf B_MIREQUESTRAMREADDATA134 (MIREQUESTRAMREADDATA_IN[134], MIREQUESTRAMREADDATA[134]);
  buf B_MIREQUESTRAMREADDATA135 (MIREQUESTRAMREADDATA_IN[135], MIREQUESTRAMREADDATA[135]);
  buf B_MIREQUESTRAMREADDATA136 (MIREQUESTRAMREADDATA_IN[136], MIREQUESTRAMREADDATA[136]);
  buf B_MIREQUESTRAMREADDATA137 (MIREQUESTRAMREADDATA_IN[137], MIREQUESTRAMREADDATA[137]);
  buf B_MIREQUESTRAMREADDATA138 (MIREQUESTRAMREADDATA_IN[138], MIREQUESTRAMREADDATA[138]);
  buf B_MIREQUESTRAMREADDATA139 (MIREQUESTRAMREADDATA_IN[139], MIREQUESTRAMREADDATA[139]);
  buf B_MIREQUESTRAMREADDATA14 (MIREQUESTRAMREADDATA_IN[14], MIREQUESTRAMREADDATA[14]);
  buf B_MIREQUESTRAMREADDATA140 (MIREQUESTRAMREADDATA_IN[140], MIREQUESTRAMREADDATA[140]);
  buf B_MIREQUESTRAMREADDATA141 (MIREQUESTRAMREADDATA_IN[141], MIREQUESTRAMREADDATA[141]);
  buf B_MIREQUESTRAMREADDATA142 (MIREQUESTRAMREADDATA_IN[142], MIREQUESTRAMREADDATA[142]);
  buf B_MIREQUESTRAMREADDATA143 (MIREQUESTRAMREADDATA_IN[143], MIREQUESTRAMREADDATA[143]);
  buf B_MIREQUESTRAMREADDATA15 (MIREQUESTRAMREADDATA_IN[15], MIREQUESTRAMREADDATA[15]);
  buf B_MIREQUESTRAMREADDATA16 (MIREQUESTRAMREADDATA_IN[16], MIREQUESTRAMREADDATA[16]);
  buf B_MIREQUESTRAMREADDATA17 (MIREQUESTRAMREADDATA_IN[17], MIREQUESTRAMREADDATA[17]);
  buf B_MIREQUESTRAMREADDATA18 (MIREQUESTRAMREADDATA_IN[18], MIREQUESTRAMREADDATA[18]);
  buf B_MIREQUESTRAMREADDATA19 (MIREQUESTRAMREADDATA_IN[19], MIREQUESTRAMREADDATA[19]);
  buf B_MIREQUESTRAMREADDATA2 (MIREQUESTRAMREADDATA_IN[2], MIREQUESTRAMREADDATA[2]);
  buf B_MIREQUESTRAMREADDATA20 (MIREQUESTRAMREADDATA_IN[20], MIREQUESTRAMREADDATA[20]);
  buf B_MIREQUESTRAMREADDATA21 (MIREQUESTRAMREADDATA_IN[21], MIREQUESTRAMREADDATA[21]);
  buf B_MIREQUESTRAMREADDATA22 (MIREQUESTRAMREADDATA_IN[22], MIREQUESTRAMREADDATA[22]);
  buf B_MIREQUESTRAMREADDATA23 (MIREQUESTRAMREADDATA_IN[23], MIREQUESTRAMREADDATA[23]);
  buf B_MIREQUESTRAMREADDATA24 (MIREQUESTRAMREADDATA_IN[24], MIREQUESTRAMREADDATA[24]);
  buf B_MIREQUESTRAMREADDATA25 (MIREQUESTRAMREADDATA_IN[25], MIREQUESTRAMREADDATA[25]);
  buf B_MIREQUESTRAMREADDATA26 (MIREQUESTRAMREADDATA_IN[26], MIREQUESTRAMREADDATA[26]);
  buf B_MIREQUESTRAMREADDATA27 (MIREQUESTRAMREADDATA_IN[27], MIREQUESTRAMREADDATA[27]);
  buf B_MIREQUESTRAMREADDATA28 (MIREQUESTRAMREADDATA_IN[28], MIREQUESTRAMREADDATA[28]);
  buf B_MIREQUESTRAMREADDATA29 (MIREQUESTRAMREADDATA_IN[29], MIREQUESTRAMREADDATA[29]);
  buf B_MIREQUESTRAMREADDATA3 (MIREQUESTRAMREADDATA_IN[3], MIREQUESTRAMREADDATA[3]);
  buf B_MIREQUESTRAMREADDATA30 (MIREQUESTRAMREADDATA_IN[30], MIREQUESTRAMREADDATA[30]);
  buf B_MIREQUESTRAMREADDATA31 (MIREQUESTRAMREADDATA_IN[31], MIREQUESTRAMREADDATA[31]);
  buf B_MIREQUESTRAMREADDATA32 (MIREQUESTRAMREADDATA_IN[32], MIREQUESTRAMREADDATA[32]);
  buf B_MIREQUESTRAMREADDATA33 (MIREQUESTRAMREADDATA_IN[33], MIREQUESTRAMREADDATA[33]);
  buf B_MIREQUESTRAMREADDATA34 (MIREQUESTRAMREADDATA_IN[34], MIREQUESTRAMREADDATA[34]);
  buf B_MIREQUESTRAMREADDATA35 (MIREQUESTRAMREADDATA_IN[35], MIREQUESTRAMREADDATA[35]);
  buf B_MIREQUESTRAMREADDATA36 (MIREQUESTRAMREADDATA_IN[36], MIREQUESTRAMREADDATA[36]);
  buf B_MIREQUESTRAMREADDATA37 (MIREQUESTRAMREADDATA_IN[37], MIREQUESTRAMREADDATA[37]);
  buf B_MIREQUESTRAMREADDATA38 (MIREQUESTRAMREADDATA_IN[38], MIREQUESTRAMREADDATA[38]);
  buf B_MIREQUESTRAMREADDATA39 (MIREQUESTRAMREADDATA_IN[39], MIREQUESTRAMREADDATA[39]);
  buf B_MIREQUESTRAMREADDATA4 (MIREQUESTRAMREADDATA_IN[4], MIREQUESTRAMREADDATA[4]);
  buf B_MIREQUESTRAMREADDATA40 (MIREQUESTRAMREADDATA_IN[40], MIREQUESTRAMREADDATA[40]);
  buf B_MIREQUESTRAMREADDATA41 (MIREQUESTRAMREADDATA_IN[41], MIREQUESTRAMREADDATA[41]);
  buf B_MIREQUESTRAMREADDATA42 (MIREQUESTRAMREADDATA_IN[42], MIREQUESTRAMREADDATA[42]);
  buf B_MIREQUESTRAMREADDATA43 (MIREQUESTRAMREADDATA_IN[43], MIREQUESTRAMREADDATA[43]);
  buf B_MIREQUESTRAMREADDATA44 (MIREQUESTRAMREADDATA_IN[44], MIREQUESTRAMREADDATA[44]);
  buf B_MIREQUESTRAMREADDATA45 (MIREQUESTRAMREADDATA_IN[45], MIREQUESTRAMREADDATA[45]);
  buf B_MIREQUESTRAMREADDATA46 (MIREQUESTRAMREADDATA_IN[46], MIREQUESTRAMREADDATA[46]);
  buf B_MIREQUESTRAMREADDATA47 (MIREQUESTRAMREADDATA_IN[47], MIREQUESTRAMREADDATA[47]);
  buf B_MIREQUESTRAMREADDATA48 (MIREQUESTRAMREADDATA_IN[48], MIREQUESTRAMREADDATA[48]);
  buf B_MIREQUESTRAMREADDATA49 (MIREQUESTRAMREADDATA_IN[49], MIREQUESTRAMREADDATA[49]);
  buf B_MIREQUESTRAMREADDATA5 (MIREQUESTRAMREADDATA_IN[5], MIREQUESTRAMREADDATA[5]);
  buf B_MIREQUESTRAMREADDATA50 (MIREQUESTRAMREADDATA_IN[50], MIREQUESTRAMREADDATA[50]);
  buf B_MIREQUESTRAMREADDATA51 (MIREQUESTRAMREADDATA_IN[51], MIREQUESTRAMREADDATA[51]);
  buf B_MIREQUESTRAMREADDATA52 (MIREQUESTRAMREADDATA_IN[52], MIREQUESTRAMREADDATA[52]);
  buf B_MIREQUESTRAMREADDATA53 (MIREQUESTRAMREADDATA_IN[53], MIREQUESTRAMREADDATA[53]);
  buf B_MIREQUESTRAMREADDATA54 (MIREQUESTRAMREADDATA_IN[54], MIREQUESTRAMREADDATA[54]);
  buf B_MIREQUESTRAMREADDATA55 (MIREQUESTRAMREADDATA_IN[55], MIREQUESTRAMREADDATA[55]);
  buf B_MIREQUESTRAMREADDATA56 (MIREQUESTRAMREADDATA_IN[56], MIREQUESTRAMREADDATA[56]);
  buf B_MIREQUESTRAMREADDATA57 (MIREQUESTRAMREADDATA_IN[57], MIREQUESTRAMREADDATA[57]);
  buf B_MIREQUESTRAMREADDATA58 (MIREQUESTRAMREADDATA_IN[58], MIREQUESTRAMREADDATA[58]);
  buf B_MIREQUESTRAMREADDATA59 (MIREQUESTRAMREADDATA_IN[59], MIREQUESTRAMREADDATA[59]);
  buf B_MIREQUESTRAMREADDATA6 (MIREQUESTRAMREADDATA_IN[6], MIREQUESTRAMREADDATA[6]);
  buf B_MIREQUESTRAMREADDATA60 (MIREQUESTRAMREADDATA_IN[60], MIREQUESTRAMREADDATA[60]);
  buf B_MIREQUESTRAMREADDATA61 (MIREQUESTRAMREADDATA_IN[61], MIREQUESTRAMREADDATA[61]);
  buf B_MIREQUESTRAMREADDATA62 (MIREQUESTRAMREADDATA_IN[62], MIREQUESTRAMREADDATA[62]);
  buf B_MIREQUESTRAMREADDATA63 (MIREQUESTRAMREADDATA_IN[63], MIREQUESTRAMREADDATA[63]);
  buf B_MIREQUESTRAMREADDATA64 (MIREQUESTRAMREADDATA_IN[64], MIREQUESTRAMREADDATA[64]);
  buf B_MIREQUESTRAMREADDATA65 (MIREQUESTRAMREADDATA_IN[65], MIREQUESTRAMREADDATA[65]);
  buf B_MIREQUESTRAMREADDATA66 (MIREQUESTRAMREADDATA_IN[66], MIREQUESTRAMREADDATA[66]);
  buf B_MIREQUESTRAMREADDATA67 (MIREQUESTRAMREADDATA_IN[67], MIREQUESTRAMREADDATA[67]);
  buf B_MIREQUESTRAMREADDATA68 (MIREQUESTRAMREADDATA_IN[68], MIREQUESTRAMREADDATA[68]);
  buf B_MIREQUESTRAMREADDATA69 (MIREQUESTRAMREADDATA_IN[69], MIREQUESTRAMREADDATA[69]);
  buf B_MIREQUESTRAMREADDATA7 (MIREQUESTRAMREADDATA_IN[7], MIREQUESTRAMREADDATA[7]);
  buf B_MIREQUESTRAMREADDATA70 (MIREQUESTRAMREADDATA_IN[70], MIREQUESTRAMREADDATA[70]);
  buf B_MIREQUESTRAMREADDATA71 (MIREQUESTRAMREADDATA_IN[71], MIREQUESTRAMREADDATA[71]);
  buf B_MIREQUESTRAMREADDATA72 (MIREQUESTRAMREADDATA_IN[72], MIREQUESTRAMREADDATA[72]);
  buf B_MIREQUESTRAMREADDATA73 (MIREQUESTRAMREADDATA_IN[73], MIREQUESTRAMREADDATA[73]);
  buf B_MIREQUESTRAMREADDATA74 (MIREQUESTRAMREADDATA_IN[74], MIREQUESTRAMREADDATA[74]);
  buf B_MIREQUESTRAMREADDATA75 (MIREQUESTRAMREADDATA_IN[75], MIREQUESTRAMREADDATA[75]);
  buf B_MIREQUESTRAMREADDATA76 (MIREQUESTRAMREADDATA_IN[76], MIREQUESTRAMREADDATA[76]);
  buf B_MIREQUESTRAMREADDATA77 (MIREQUESTRAMREADDATA_IN[77], MIREQUESTRAMREADDATA[77]);
  buf B_MIREQUESTRAMREADDATA78 (MIREQUESTRAMREADDATA_IN[78], MIREQUESTRAMREADDATA[78]);
  buf B_MIREQUESTRAMREADDATA79 (MIREQUESTRAMREADDATA_IN[79], MIREQUESTRAMREADDATA[79]);
  buf B_MIREQUESTRAMREADDATA8 (MIREQUESTRAMREADDATA_IN[8], MIREQUESTRAMREADDATA[8]);
  buf B_MIREQUESTRAMREADDATA80 (MIREQUESTRAMREADDATA_IN[80], MIREQUESTRAMREADDATA[80]);
  buf B_MIREQUESTRAMREADDATA81 (MIREQUESTRAMREADDATA_IN[81], MIREQUESTRAMREADDATA[81]);
  buf B_MIREQUESTRAMREADDATA82 (MIREQUESTRAMREADDATA_IN[82], MIREQUESTRAMREADDATA[82]);
  buf B_MIREQUESTRAMREADDATA83 (MIREQUESTRAMREADDATA_IN[83], MIREQUESTRAMREADDATA[83]);
  buf B_MIREQUESTRAMREADDATA84 (MIREQUESTRAMREADDATA_IN[84], MIREQUESTRAMREADDATA[84]);
  buf B_MIREQUESTRAMREADDATA85 (MIREQUESTRAMREADDATA_IN[85], MIREQUESTRAMREADDATA[85]);
  buf B_MIREQUESTRAMREADDATA86 (MIREQUESTRAMREADDATA_IN[86], MIREQUESTRAMREADDATA[86]);
  buf B_MIREQUESTRAMREADDATA87 (MIREQUESTRAMREADDATA_IN[87], MIREQUESTRAMREADDATA[87]);
  buf B_MIREQUESTRAMREADDATA88 (MIREQUESTRAMREADDATA_IN[88], MIREQUESTRAMREADDATA[88]);
  buf B_MIREQUESTRAMREADDATA89 (MIREQUESTRAMREADDATA_IN[89], MIREQUESTRAMREADDATA[89]);
  buf B_MIREQUESTRAMREADDATA9 (MIREQUESTRAMREADDATA_IN[9], MIREQUESTRAMREADDATA[9]);
  buf B_MIREQUESTRAMREADDATA90 (MIREQUESTRAMREADDATA_IN[90], MIREQUESTRAMREADDATA[90]);
  buf B_MIREQUESTRAMREADDATA91 (MIREQUESTRAMREADDATA_IN[91], MIREQUESTRAMREADDATA[91]);
  buf B_MIREQUESTRAMREADDATA92 (MIREQUESTRAMREADDATA_IN[92], MIREQUESTRAMREADDATA[92]);
  buf B_MIREQUESTRAMREADDATA93 (MIREQUESTRAMREADDATA_IN[93], MIREQUESTRAMREADDATA[93]);
  buf B_MIREQUESTRAMREADDATA94 (MIREQUESTRAMREADDATA_IN[94], MIREQUESTRAMREADDATA[94]);
  buf B_MIREQUESTRAMREADDATA95 (MIREQUESTRAMREADDATA_IN[95], MIREQUESTRAMREADDATA[95]);
  buf B_MIREQUESTRAMREADDATA96 (MIREQUESTRAMREADDATA_IN[96], MIREQUESTRAMREADDATA[96]);
  buf B_MIREQUESTRAMREADDATA97 (MIREQUESTRAMREADDATA_IN[97], MIREQUESTRAMREADDATA[97]);
  buf B_MIREQUESTRAMREADDATA98 (MIREQUESTRAMREADDATA_IN[98], MIREQUESTRAMREADDATA[98]);
  buf B_MIREQUESTRAMREADDATA99 (MIREQUESTRAMREADDATA_IN[99], MIREQUESTRAMREADDATA[99]);
  buf B_PCIECQNPREQ (PCIECQNPREQ_IN, PCIECQNPREQ);
  buf B_PIPECLK (PIPECLK_IN, PIPECLK);
  buf B_PIPEEQFS0 (PIPEEQFS_IN[0], PIPEEQFS[0]);
  buf B_PIPEEQFS1 (PIPEEQFS_IN[1], PIPEEQFS[1]);
  buf B_PIPEEQFS2 (PIPEEQFS_IN[2], PIPEEQFS[2]);
  buf B_PIPEEQFS3 (PIPEEQFS_IN[3], PIPEEQFS[3]);
  buf B_PIPEEQFS4 (PIPEEQFS_IN[4], PIPEEQFS[4]);
  buf B_PIPEEQFS5 (PIPEEQFS_IN[5], PIPEEQFS[5]);
  buf B_PIPEEQLF0 (PIPEEQLF_IN[0], PIPEEQLF[0]);
  buf B_PIPEEQLF1 (PIPEEQLF_IN[1], PIPEEQLF[1]);
  buf B_PIPEEQLF2 (PIPEEQLF_IN[2], PIPEEQLF[2]);
  buf B_PIPEEQLF3 (PIPEEQLF_IN[3], PIPEEQLF[3]);
  buf B_PIPEEQLF4 (PIPEEQLF_IN[4], PIPEEQLF[4]);
  buf B_PIPEEQLF5 (PIPEEQLF_IN[5], PIPEEQLF[5]);
  buf B_PIPERESETN (PIPERESETN_IN, PIPERESETN);
  buf B_PIPERX0CHARISK0 (PIPERX0CHARISK_IN[0], PIPERX0CHARISK[0]);
  buf B_PIPERX0CHARISK1 (PIPERX0CHARISK_IN[1], PIPERX0CHARISK[1]);
  buf B_PIPERX0DATA0 (PIPERX0DATA_IN[0], PIPERX0DATA[0]);
  buf B_PIPERX0DATA1 (PIPERX0DATA_IN[1], PIPERX0DATA[1]);
  buf B_PIPERX0DATA10 (PIPERX0DATA_IN[10], PIPERX0DATA[10]);
  buf B_PIPERX0DATA11 (PIPERX0DATA_IN[11], PIPERX0DATA[11]);
  buf B_PIPERX0DATA12 (PIPERX0DATA_IN[12], PIPERX0DATA[12]);
  buf B_PIPERX0DATA13 (PIPERX0DATA_IN[13], PIPERX0DATA[13]);
  buf B_PIPERX0DATA14 (PIPERX0DATA_IN[14], PIPERX0DATA[14]);
  buf B_PIPERX0DATA15 (PIPERX0DATA_IN[15], PIPERX0DATA[15]);
  buf B_PIPERX0DATA16 (PIPERX0DATA_IN[16], PIPERX0DATA[16]);
  buf B_PIPERX0DATA17 (PIPERX0DATA_IN[17], PIPERX0DATA[17]);
  buf B_PIPERX0DATA18 (PIPERX0DATA_IN[18], PIPERX0DATA[18]);
  buf B_PIPERX0DATA19 (PIPERX0DATA_IN[19], PIPERX0DATA[19]);
  buf B_PIPERX0DATA2 (PIPERX0DATA_IN[2], PIPERX0DATA[2]);
  buf B_PIPERX0DATA20 (PIPERX0DATA_IN[20], PIPERX0DATA[20]);
  buf B_PIPERX0DATA21 (PIPERX0DATA_IN[21], PIPERX0DATA[21]);
  buf B_PIPERX0DATA22 (PIPERX0DATA_IN[22], PIPERX0DATA[22]);
  buf B_PIPERX0DATA23 (PIPERX0DATA_IN[23], PIPERX0DATA[23]);
  buf B_PIPERX0DATA24 (PIPERX0DATA_IN[24], PIPERX0DATA[24]);
  buf B_PIPERX0DATA25 (PIPERX0DATA_IN[25], PIPERX0DATA[25]);
  buf B_PIPERX0DATA26 (PIPERX0DATA_IN[26], PIPERX0DATA[26]);
  buf B_PIPERX0DATA27 (PIPERX0DATA_IN[27], PIPERX0DATA[27]);
  buf B_PIPERX0DATA28 (PIPERX0DATA_IN[28], PIPERX0DATA[28]);
  buf B_PIPERX0DATA29 (PIPERX0DATA_IN[29], PIPERX0DATA[29]);
  buf B_PIPERX0DATA3 (PIPERX0DATA_IN[3], PIPERX0DATA[3]);
  buf B_PIPERX0DATA30 (PIPERX0DATA_IN[30], PIPERX0DATA[30]);
  buf B_PIPERX0DATA31 (PIPERX0DATA_IN[31], PIPERX0DATA[31]);
  buf B_PIPERX0DATA4 (PIPERX0DATA_IN[4], PIPERX0DATA[4]);
  buf B_PIPERX0DATA5 (PIPERX0DATA_IN[5], PIPERX0DATA[5]);
  buf B_PIPERX0DATA6 (PIPERX0DATA_IN[6], PIPERX0DATA[6]);
  buf B_PIPERX0DATA7 (PIPERX0DATA_IN[7], PIPERX0DATA[7]);
  buf B_PIPERX0DATA8 (PIPERX0DATA_IN[8], PIPERX0DATA[8]);
  buf B_PIPERX0DATA9 (PIPERX0DATA_IN[9], PIPERX0DATA[9]);
  buf B_PIPERX0DATAVALID (PIPERX0DATAVALID_IN, PIPERX0DATAVALID);
  buf B_PIPERX0ELECIDLE (PIPERX0ELECIDLE_IN, PIPERX0ELECIDLE);
  buf B_PIPERX0EQDONE (PIPERX0EQDONE_IN, PIPERX0EQDONE);
  buf B_PIPERX0EQLPADAPTDONE (PIPERX0EQLPADAPTDONE_IN, PIPERX0EQLPADAPTDONE);
  buf B_PIPERX0EQLPLFFSSEL (PIPERX0EQLPLFFSSEL_IN, PIPERX0EQLPLFFSSEL);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET0 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[0], PIPERX0EQLPNEWTXCOEFFORPRESET[0]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET1 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[1], PIPERX0EQLPNEWTXCOEFFORPRESET[1]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET10 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[10], PIPERX0EQLPNEWTXCOEFFORPRESET[10]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET11 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[11], PIPERX0EQLPNEWTXCOEFFORPRESET[11]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET12 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[12], PIPERX0EQLPNEWTXCOEFFORPRESET[12]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET13 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[13], PIPERX0EQLPNEWTXCOEFFORPRESET[13]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET14 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[14], PIPERX0EQLPNEWTXCOEFFORPRESET[14]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET15 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[15], PIPERX0EQLPNEWTXCOEFFORPRESET[15]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET16 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[16], PIPERX0EQLPNEWTXCOEFFORPRESET[16]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET17 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[17], PIPERX0EQLPNEWTXCOEFFORPRESET[17]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET2 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[2], PIPERX0EQLPNEWTXCOEFFORPRESET[2]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET3 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[3], PIPERX0EQLPNEWTXCOEFFORPRESET[3]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET4 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[4], PIPERX0EQLPNEWTXCOEFFORPRESET[4]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET5 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[5], PIPERX0EQLPNEWTXCOEFFORPRESET[5]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET6 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[6], PIPERX0EQLPNEWTXCOEFFORPRESET[6]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET7 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[7], PIPERX0EQLPNEWTXCOEFFORPRESET[7]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET8 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[8], PIPERX0EQLPNEWTXCOEFFORPRESET[8]);
  buf B_PIPERX0EQLPNEWTXCOEFFORPRESET9 (PIPERX0EQLPNEWTXCOEFFORPRESET_IN[9], PIPERX0EQLPNEWTXCOEFFORPRESET[9]);
  buf B_PIPERX0PHYSTATUS (PIPERX0PHYSTATUS_IN, PIPERX0PHYSTATUS);
  buf B_PIPERX0STARTBLOCK (PIPERX0STARTBLOCK_IN, PIPERX0STARTBLOCK);
  buf B_PIPERX0STATUS0 (PIPERX0STATUS_IN[0], PIPERX0STATUS[0]);
  buf B_PIPERX0STATUS1 (PIPERX0STATUS_IN[1], PIPERX0STATUS[1]);
  buf B_PIPERX0STATUS2 (PIPERX0STATUS_IN[2], PIPERX0STATUS[2]);
  buf B_PIPERX0SYNCHEADER0 (PIPERX0SYNCHEADER_IN[0], PIPERX0SYNCHEADER[0]);
  buf B_PIPERX0SYNCHEADER1 (PIPERX0SYNCHEADER_IN[1], PIPERX0SYNCHEADER[1]);
  buf B_PIPERX0VALID (PIPERX0VALID_IN, PIPERX0VALID);
  buf B_PIPERX1CHARISK0 (PIPERX1CHARISK_IN[0], PIPERX1CHARISK[0]);
  buf B_PIPERX1CHARISK1 (PIPERX1CHARISK_IN[1], PIPERX1CHARISK[1]);
  buf B_PIPERX1DATA0 (PIPERX1DATA_IN[0], PIPERX1DATA[0]);
  buf B_PIPERX1DATA1 (PIPERX1DATA_IN[1], PIPERX1DATA[1]);
  buf B_PIPERX1DATA10 (PIPERX1DATA_IN[10], PIPERX1DATA[10]);
  buf B_PIPERX1DATA11 (PIPERX1DATA_IN[11], PIPERX1DATA[11]);
  buf B_PIPERX1DATA12 (PIPERX1DATA_IN[12], PIPERX1DATA[12]);
  buf B_PIPERX1DATA13 (PIPERX1DATA_IN[13], PIPERX1DATA[13]);
  buf B_PIPERX1DATA14 (PIPERX1DATA_IN[14], PIPERX1DATA[14]);
  buf B_PIPERX1DATA15 (PIPERX1DATA_IN[15], PIPERX1DATA[15]);
  buf B_PIPERX1DATA16 (PIPERX1DATA_IN[16], PIPERX1DATA[16]);
  buf B_PIPERX1DATA17 (PIPERX1DATA_IN[17], PIPERX1DATA[17]);
  buf B_PIPERX1DATA18 (PIPERX1DATA_IN[18], PIPERX1DATA[18]);
  buf B_PIPERX1DATA19 (PIPERX1DATA_IN[19], PIPERX1DATA[19]);
  buf B_PIPERX1DATA2 (PIPERX1DATA_IN[2], PIPERX1DATA[2]);
  buf B_PIPERX1DATA20 (PIPERX1DATA_IN[20], PIPERX1DATA[20]);
  buf B_PIPERX1DATA21 (PIPERX1DATA_IN[21], PIPERX1DATA[21]);
  buf B_PIPERX1DATA22 (PIPERX1DATA_IN[22], PIPERX1DATA[22]);
  buf B_PIPERX1DATA23 (PIPERX1DATA_IN[23], PIPERX1DATA[23]);
  buf B_PIPERX1DATA24 (PIPERX1DATA_IN[24], PIPERX1DATA[24]);
  buf B_PIPERX1DATA25 (PIPERX1DATA_IN[25], PIPERX1DATA[25]);
  buf B_PIPERX1DATA26 (PIPERX1DATA_IN[26], PIPERX1DATA[26]);
  buf B_PIPERX1DATA27 (PIPERX1DATA_IN[27], PIPERX1DATA[27]);
  buf B_PIPERX1DATA28 (PIPERX1DATA_IN[28], PIPERX1DATA[28]);
  buf B_PIPERX1DATA29 (PIPERX1DATA_IN[29], PIPERX1DATA[29]);
  buf B_PIPERX1DATA3 (PIPERX1DATA_IN[3], PIPERX1DATA[3]);
  buf B_PIPERX1DATA30 (PIPERX1DATA_IN[30], PIPERX1DATA[30]);
  buf B_PIPERX1DATA31 (PIPERX1DATA_IN[31], PIPERX1DATA[31]);
  buf B_PIPERX1DATA4 (PIPERX1DATA_IN[4], PIPERX1DATA[4]);
  buf B_PIPERX1DATA5 (PIPERX1DATA_IN[5], PIPERX1DATA[5]);
  buf B_PIPERX1DATA6 (PIPERX1DATA_IN[6], PIPERX1DATA[6]);
  buf B_PIPERX1DATA7 (PIPERX1DATA_IN[7], PIPERX1DATA[7]);
  buf B_PIPERX1DATA8 (PIPERX1DATA_IN[8], PIPERX1DATA[8]);
  buf B_PIPERX1DATA9 (PIPERX1DATA_IN[9], PIPERX1DATA[9]);
  buf B_PIPERX1DATAVALID (PIPERX1DATAVALID_IN, PIPERX1DATAVALID);
  buf B_PIPERX1ELECIDLE (PIPERX1ELECIDLE_IN, PIPERX1ELECIDLE);
  buf B_PIPERX1EQDONE (PIPERX1EQDONE_IN, PIPERX1EQDONE);
  buf B_PIPERX1EQLPADAPTDONE (PIPERX1EQLPADAPTDONE_IN, PIPERX1EQLPADAPTDONE);
  buf B_PIPERX1EQLPLFFSSEL (PIPERX1EQLPLFFSSEL_IN, PIPERX1EQLPLFFSSEL);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET0 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[0], PIPERX1EQLPNEWTXCOEFFORPRESET[0]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET1 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[1], PIPERX1EQLPNEWTXCOEFFORPRESET[1]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET10 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[10], PIPERX1EQLPNEWTXCOEFFORPRESET[10]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET11 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[11], PIPERX1EQLPNEWTXCOEFFORPRESET[11]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET12 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[12], PIPERX1EQLPNEWTXCOEFFORPRESET[12]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET13 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[13], PIPERX1EQLPNEWTXCOEFFORPRESET[13]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET14 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[14], PIPERX1EQLPNEWTXCOEFFORPRESET[14]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET15 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[15], PIPERX1EQLPNEWTXCOEFFORPRESET[15]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET16 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[16], PIPERX1EQLPNEWTXCOEFFORPRESET[16]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET17 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[17], PIPERX1EQLPNEWTXCOEFFORPRESET[17]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET2 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[2], PIPERX1EQLPNEWTXCOEFFORPRESET[2]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET3 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[3], PIPERX1EQLPNEWTXCOEFFORPRESET[3]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET4 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[4], PIPERX1EQLPNEWTXCOEFFORPRESET[4]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET5 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[5], PIPERX1EQLPNEWTXCOEFFORPRESET[5]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET6 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[6], PIPERX1EQLPNEWTXCOEFFORPRESET[6]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET7 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[7], PIPERX1EQLPNEWTXCOEFFORPRESET[7]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET8 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[8], PIPERX1EQLPNEWTXCOEFFORPRESET[8]);
  buf B_PIPERX1EQLPNEWTXCOEFFORPRESET9 (PIPERX1EQLPNEWTXCOEFFORPRESET_IN[9], PIPERX1EQLPNEWTXCOEFFORPRESET[9]);
  buf B_PIPERX1PHYSTATUS (PIPERX1PHYSTATUS_IN, PIPERX1PHYSTATUS);
  buf B_PIPERX1STARTBLOCK (PIPERX1STARTBLOCK_IN, PIPERX1STARTBLOCK);
  buf B_PIPERX1STATUS0 (PIPERX1STATUS_IN[0], PIPERX1STATUS[0]);
  buf B_PIPERX1STATUS1 (PIPERX1STATUS_IN[1], PIPERX1STATUS[1]);
  buf B_PIPERX1STATUS2 (PIPERX1STATUS_IN[2], PIPERX1STATUS[2]);
  buf B_PIPERX1SYNCHEADER0 (PIPERX1SYNCHEADER_IN[0], PIPERX1SYNCHEADER[0]);
  buf B_PIPERX1SYNCHEADER1 (PIPERX1SYNCHEADER_IN[1], PIPERX1SYNCHEADER[1]);
  buf B_PIPERX1VALID (PIPERX1VALID_IN, PIPERX1VALID);
  buf B_PIPERX2CHARISK0 (PIPERX2CHARISK_IN[0], PIPERX2CHARISK[0]);
  buf B_PIPERX2CHARISK1 (PIPERX2CHARISK_IN[1], PIPERX2CHARISK[1]);
  buf B_PIPERX2DATA0 (PIPERX2DATA_IN[0], PIPERX2DATA[0]);
  buf B_PIPERX2DATA1 (PIPERX2DATA_IN[1], PIPERX2DATA[1]);
  buf B_PIPERX2DATA10 (PIPERX2DATA_IN[10], PIPERX2DATA[10]);
  buf B_PIPERX2DATA11 (PIPERX2DATA_IN[11], PIPERX2DATA[11]);
  buf B_PIPERX2DATA12 (PIPERX2DATA_IN[12], PIPERX2DATA[12]);
  buf B_PIPERX2DATA13 (PIPERX2DATA_IN[13], PIPERX2DATA[13]);
  buf B_PIPERX2DATA14 (PIPERX2DATA_IN[14], PIPERX2DATA[14]);
  buf B_PIPERX2DATA15 (PIPERX2DATA_IN[15], PIPERX2DATA[15]);
  buf B_PIPERX2DATA16 (PIPERX2DATA_IN[16], PIPERX2DATA[16]);
  buf B_PIPERX2DATA17 (PIPERX2DATA_IN[17], PIPERX2DATA[17]);
  buf B_PIPERX2DATA18 (PIPERX2DATA_IN[18], PIPERX2DATA[18]);
  buf B_PIPERX2DATA19 (PIPERX2DATA_IN[19], PIPERX2DATA[19]);
  buf B_PIPERX2DATA2 (PIPERX2DATA_IN[2], PIPERX2DATA[2]);
  buf B_PIPERX2DATA20 (PIPERX2DATA_IN[20], PIPERX2DATA[20]);
  buf B_PIPERX2DATA21 (PIPERX2DATA_IN[21], PIPERX2DATA[21]);
  buf B_PIPERX2DATA22 (PIPERX2DATA_IN[22], PIPERX2DATA[22]);
  buf B_PIPERX2DATA23 (PIPERX2DATA_IN[23], PIPERX2DATA[23]);
  buf B_PIPERX2DATA24 (PIPERX2DATA_IN[24], PIPERX2DATA[24]);
  buf B_PIPERX2DATA25 (PIPERX2DATA_IN[25], PIPERX2DATA[25]);
  buf B_PIPERX2DATA26 (PIPERX2DATA_IN[26], PIPERX2DATA[26]);
  buf B_PIPERX2DATA27 (PIPERX2DATA_IN[27], PIPERX2DATA[27]);
  buf B_PIPERX2DATA28 (PIPERX2DATA_IN[28], PIPERX2DATA[28]);
  buf B_PIPERX2DATA29 (PIPERX2DATA_IN[29], PIPERX2DATA[29]);
  buf B_PIPERX2DATA3 (PIPERX2DATA_IN[3], PIPERX2DATA[3]);
  buf B_PIPERX2DATA30 (PIPERX2DATA_IN[30], PIPERX2DATA[30]);
  buf B_PIPERX2DATA31 (PIPERX2DATA_IN[31], PIPERX2DATA[31]);
  buf B_PIPERX2DATA4 (PIPERX2DATA_IN[4], PIPERX2DATA[4]);
  buf B_PIPERX2DATA5 (PIPERX2DATA_IN[5], PIPERX2DATA[5]);
  buf B_PIPERX2DATA6 (PIPERX2DATA_IN[6], PIPERX2DATA[6]);
  buf B_PIPERX2DATA7 (PIPERX2DATA_IN[7], PIPERX2DATA[7]);
  buf B_PIPERX2DATA8 (PIPERX2DATA_IN[8], PIPERX2DATA[8]);
  buf B_PIPERX2DATA9 (PIPERX2DATA_IN[9], PIPERX2DATA[9]);
  buf B_PIPERX2DATAVALID (PIPERX2DATAVALID_IN, PIPERX2DATAVALID);
  buf B_PIPERX2ELECIDLE (PIPERX2ELECIDLE_IN, PIPERX2ELECIDLE);
  buf B_PIPERX2EQDONE (PIPERX2EQDONE_IN, PIPERX2EQDONE);
  buf B_PIPERX2EQLPADAPTDONE (PIPERX2EQLPADAPTDONE_IN, PIPERX2EQLPADAPTDONE);
  buf B_PIPERX2EQLPLFFSSEL (PIPERX2EQLPLFFSSEL_IN, PIPERX2EQLPLFFSSEL);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET0 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[0], PIPERX2EQLPNEWTXCOEFFORPRESET[0]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET1 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[1], PIPERX2EQLPNEWTXCOEFFORPRESET[1]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET10 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[10], PIPERX2EQLPNEWTXCOEFFORPRESET[10]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET11 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[11], PIPERX2EQLPNEWTXCOEFFORPRESET[11]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET12 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[12], PIPERX2EQLPNEWTXCOEFFORPRESET[12]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET13 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[13], PIPERX2EQLPNEWTXCOEFFORPRESET[13]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET14 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[14], PIPERX2EQLPNEWTXCOEFFORPRESET[14]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET15 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[15], PIPERX2EQLPNEWTXCOEFFORPRESET[15]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET16 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[16], PIPERX2EQLPNEWTXCOEFFORPRESET[16]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET17 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[17], PIPERX2EQLPNEWTXCOEFFORPRESET[17]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET2 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[2], PIPERX2EQLPNEWTXCOEFFORPRESET[2]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET3 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[3], PIPERX2EQLPNEWTXCOEFFORPRESET[3]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET4 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[4], PIPERX2EQLPNEWTXCOEFFORPRESET[4]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET5 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[5], PIPERX2EQLPNEWTXCOEFFORPRESET[5]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET6 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[6], PIPERX2EQLPNEWTXCOEFFORPRESET[6]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET7 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[7], PIPERX2EQLPNEWTXCOEFFORPRESET[7]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET8 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[8], PIPERX2EQLPNEWTXCOEFFORPRESET[8]);
  buf B_PIPERX2EQLPNEWTXCOEFFORPRESET9 (PIPERX2EQLPNEWTXCOEFFORPRESET_IN[9], PIPERX2EQLPNEWTXCOEFFORPRESET[9]);
  buf B_PIPERX2PHYSTATUS (PIPERX2PHYSTATUS_IN, PIPERX2PHYSTATUS);
  buf B_PIPERX2STARTBLOCK (PIPERX2STARTBLOCK_IN, PIPERX2STARTBLOCK);
  buf B_PIPERX2STATUS0 (PIPERX2STATUS_IN[0], PIPERX2STATUS[0]);
  buf B_PIPERX2STATUS1 (PIPERX2STATUS_IN[1], PIPERX2STATUS[1]);
  buf B_PIPERX2STATUS2 (PIPERX2STATUS_IN[2], PIPERX2STATUS[2]);
  buf B_PIPERX2SYNCHEADER0 (PIPERX2SYNCHEADER_IN[0], PIPERX2SYNCHEADER[0]);
  buf B_PIPERX2SYNCHEADER1 (PIPERX2SYNCHEADER_IN[1], PIPERX2SYNCHEADER[1]);
  buf B_PIPERX2VALID (PIPERX2VALID_IN, PIPERX2VALID);
  buf B_PIPERX3CHARISK0 (PIPERX3CHARISK_IN[0], PIPERX3CHARISK[0]);
  buf B_PIPERX3CHARISK1 (PIPERX3CHARISK_IN[1], PIPERX3CHARISK[1]);
  buf B_PIPERX3DATA0 (PIPERX3DATA_IN[0], PIPERX3DATA[0]);
  buf B_PIPERX3DATA1 (PIPERX3DATA_IN[1], PIPERX3DATA[1]);
  buf B_PIPERX3DATA10 (PIPERX3DATA_IN[10], PIPERX3DATA[10]);
  buf B_PIPERX3DATA11 (PIPERX3DATA_IN[11], PIPERX3DATA[11]);
  buf B_PIPERX3DATA12 (PIPERX3DATA_IN[12], PIPERX3DATA[12]);
  buf B_PIPERX3DATA13 (PIPERX3DATA_IN[13], PIPERX3DATA[13]);
  buf B_PIPERX3DATA14 (PIPERX3DATA_IN[14], PIPERX3DATA[14]);
  buf B_PIPERX3DATA15 (PIPERX3DATA_IN[15], PIPERX3DATA[15]);
  buf B_PIPERX3DATA16 (PIPERX3DATA_IN[16], PIPERX3DATA[16]);
  buf B_PIPERX3DATA17 (PIPERX3DATA_IN[17], PIPERX3DATA[17]);
  buf B_PIPERX3DATA18 (PIPERX3DATA_IN[18], PIPERX3DATA[18]);
  buf B_PIPERX3DATA19 (PIPERX3DATA_IN[19], PIPERX3DATA[19]);
  buf B_PIPERX3DATA2 (PIPERX3DATA_IN[2], PIPERX3DATA[2]);
  buf B_PIPERX3DATA20 (PIPERX3DATA_IN[20], PIPERX3DATA[20]);
  buf B_PIPERX3DATA21 (PIPERX3DATA_IN[21], PIPERX3DATA[21]);
  buf B_PIPERX3DATA22 (PIPERX3DATA_IN[22], PIPERX3DATA[22]);
  buf B_PIPERX3DATA23 (PIPERX3DATA_IN[23], PIPERX3DATA[23]);
  buf B_PIPERX3DATA24 (PIPERX3DATA_IN[24], PIPERX3DATA[24]);
  buf B_PIPERX3DATA25 (PIPERX3DATA_IN[25], PIPERX3DATA[25]);
  buf B_PIPERX3DATA26 (PIPERX3DATA_IN[26], PIPERX3DATA[26]);
  buf B_PIPERX3DATA27 (PIPERX3DATA_IN[27], PIPERX3DATA[27]);
  buf B_PIPERX3DATA28 (PIPERX3DATA_IN[28], PIPERX3DATA[28]);
  buf B_PIPERX3DATA29 (PIPERX3DATA_IN[29], PIPERX3DATA[29]);
  buf B_PIPERX3DATA3 (PIPERX3DATA_IN[3], PIPERX3DATA[3]);
  buf B_PIPERX3DATA30 (PIPERX3DATA_IN[30], PIPERX3DATA[30]);
  buf B_PIPERX3DATA31 (PIPERX3DATA_IN[31], PIPERX3DATA[31]);
  buf B_PIPERX3DATA4 (PIPERX3DATA_IN[4], PIPERX3DATA[4]);
  buf B_PIPERX3DATA5 (PIPERX3DATA_IN[5], PIPERX3DATA[5]);
  buf B_PIPERX3DATA6 (PIPERX3DATA_IN[6], PIPERX3DATA[6]);
  buf B_PIPERX3DATA7 (PIPERX3DATA_IN[7], PIPERX3DATA[7]);
  buf B_PIPERX3DATA8 (PIPERX3DATA_IN[8], PIPERX3DATA[8]);
  buf B_PIPERX3DATA9 (PIPERX3DATA_IN[9], PIPERX3DATA[9]);
  buf B_PIPERX3DATAVALID (PIPERX3DATAVALID_IN, PIPERX3DATAVALID);
  buf B_PIPERX3ELECIDLE (PIPERX3ELECIDLE_IN, PIPERX3ELECIDLE);
  buf B_PIPERX3EQDONE (PIPERX3EQDONE_IN, PIPERX3EQDONE);
  buf B_PIPERX3EQLPADAPTDONE (PIPERX3EQLPADAPTDONE_IN, PIPERX3EQLPADAPTDONE);
  buf B_PIPERX3EQLPLFFSSEL (PIPERX3EQLPLFFSSEL_IN, PIPERX3EQLPLFFSSEL);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET0 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[0], PIPERX3EQLPNEWTXCOEFFORPRESET[0]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET1 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[1], PIPERX3EQLPNEWTXCOEFFORPRESET[1]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET10 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[10], PIPERX3EQLPNEWTXCOEFFORPRESET[10]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET11 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[11], PIPERX3EQLPNEWTXCOEFFORPRESET[11]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET12 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[12], PIPERX3EQLPNEWTXCOEFFORPRESET[12]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET13 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[13], PIPERX3EQLPNEWTXCOEFFORPRESET[13]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET14 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[14], PIPERX3EQLPNEWTXCOEFFORPRESET[14]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET15 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[15], PIPERX3EQLPNEWTXCOEFFORPRESET[15]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET16 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[16], PIPERX3EQLPNEWTXCOEFFORPRESET[16]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET17 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[17], PIPERX3EQLPNEWTXCOEFFORPRESET[17]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET2 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[2], PIPERX3EQLPNEWTXCOEFFORPRESET[2]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET3 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[3], PIPERX3EQLPNEWTXCOEFFORPRESET[3]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET4 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[4], PIPERX3EQLPNEWTXCOEFFORPRESET[4]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET5 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[5], PIPERX3EQLPNEWTXCOEFFORPRESET[5]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET6 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[6], PIPERX3EQLPNEWTXCOEFFORPRESET[6]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET7 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[7], PIPERX3EQLPNEWTXCOEFFORPRESET[7]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET8 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[8], PIPERX3EQLPNEWTXCOEFFORPRESET[8]);
  buf B_PIPERX3EQLPNEWTXCOEFFORPRESET9 (PIPERX3EQLPNEWTXCOEFFORPRESET_IN[9], PIPERX3EQLPNEWTXCOEFFORPRESET[9]);
  buf B_PIPERX3PHYSTATUS (PIPERX3PHYSTATUS_IN, PIPERX3PHYSTATUS);
  buf B_PIPERX3STARTBLOCK (PIPERX3STARTBLOCK_IN, PIPERX3STARTBLOCK);
  buf B_PIPERX3STATUS0 (PIPERX3STATUS_IN[0], PIPERX3STATUS[0]);
  buf B_PIPERX3STATUS1 (PIPERX3STATUS_IN[1], PIPERX3STATUS[1]);
  buf B_PIPERX3STATUS2 (PIPERX3STATUS_IN[2], PIPERX3STATUS[2]);
  buf B_PIPERX3SYNCHEADER0 (PIPERX3SYNCHEADER_IN[0], PIPERX3SYNCHEADER[0]);
  buf B_PIPERX3SYNCHEADER1 (PIPERX3SYNCHEADER_IN[1], PIPERX3SYNCHEADER[1]);
  buf B_PIPERX3VALID (PIPERX3VALID_IN, PIPERX3VALID);
  buf B_PIPERX4CHARISK0 (PIPERX4CHARISK_IN[0], PIPERX4CHARISK[0]);
  buf B_PIPERX4CHARISK1 (PIPERX4CHARISK_IN[1], PIPERX4CHARISK[1]);
  buf B_PIPERX4DATA0 (PIPERX4DATA_IN[0], PIPERX4DATA[0]);
  buf B_PIPERX4DATA1 (PIPERX4DATA_IN[1], PIPERX4DATA[1]);
  buf B_PIPERX4DATA10 (PIPERX4DATA_IN[10], PIPERX4DATA[10]);
  buf B_PIPERX4DATA11 (PIPERX4DATA_IN[11], PIPERX4DATA[11]);
  buf B_PIPERX4DATA12 (PIPERX4DATA_IN[12], PIPERX4DATA[12]);
  buf B_PIPERX4DATA13 (PIPERX4DATA_IN[13], PIPERX4DATA[13]);
  buf B_PIPERX4DATA14 (PIPERX4DATA_IN[14], PIPERX4DATA[14]);
  buf B_PIPERX4DATA15 (PIPERX4DATA_IN[15], PIPERX4DATA[15]);
  buf B_PIPERX4DATA16 (PIPERX4DATA_IN[16], PIPERX4DATA[16]);
  buf B_PIPERX4DATA17 (PIPERX4DATA_IN[17], PIPERX4DATA[17]);
  buf B_PIPERX4DATA18 (PIPERX4DATA_IN[18], PIPERX4DATA[18]);
  buf B_PIPERX4DATA19 (PIPERX4DATA_IN[19], PIPERX4DATA[19]);
  buf B_PIPERX4DATA2 (PIPERX4DATA_IN[2], PIPERX4DATA[2]);
  buf B_PIPERX4DATA20 (PIPERX4DATA_IN[20], PIPERX4DATA[20]);
  buf B_PIPERX4DATA21 (PIPERX4DATA_IN[21], PIPERX4DATA[21]);
  buf B_PIPERX4DATA22 (PIPERX4DATA_IN[22], PIPERX4DATA[22]);
  buf B_PIPERX4DATA23 (PIPERX4DATA_IN[23], PIPERX4DATA[23]);
  buf B_PIPERX4DATA24 (PIPERX4DATA_IN[24], PIPERX4DATA[24]);
  buf B_PIPERX4DATA25 (PIPERX4DATA_IN[25], PIPERX4DATA[25]);
  buf B_PIPERX4DATA26 (PIPERX4DATA_IN[26], PIPERX4DATA[26]);
  buf B_PIPERX4DATA27 (PIPERX4DATA_IN[27], PIPERX4DATA[27]);
  buf B_PIPERX4DATA28 (PIPERX4DATA_IN[28], PIPERX4DATA[28]);
  buf B_PIPERX4DATA29 (PIPERX4DATA_IN[29], PIPERX4DATA[29]);
  buf B_PIPERX4DATA3 (PIPERX4DATA_IN[3], PIPERX4DATA[3]);
  buf B_PIPERX4DATA30 (PIPERX4DATA_IN[30], PIPERX4DATA[30]);
  buf B_PIPERX4DATA31 (PIPERX4DATA_IN[31], PIPERX4DATA[31]);
  buf B_PIPERX4DATA4 (PIPERX4DATA_IN[4], PIPERX4DATA[4]);
  buf B_PIPERX4DATA5 (PIPERX4DATA_IN[5], PIPERX4DATA[5]);
  buf B_PIPERX4DATA6 (PIPERX4DATA_IN[6], PIPERX4DATA[6]);
  buf B_PIPERX4DATA7 (PIPERX4DATA_IN[7], PIPERX4DATA[7]);
  buf B_PIPERX4DATA8 (PIPERX4DATA_IN[8], PIPERX4DATA[8]);
  buf B_PIPERX4DATA9 (PIPERX4DATA_IN[9], PIPERX4DATA[9]);
  buf B_PIPERX4DATAVALID (PIPERX4DATAVALID_IN, PIPERX4DATAVALID);
  buf B_PIPERX4ELECIDLE (PIPERX4ELECIDLE_IN, PIPERX4ELECIDLE);
  buf B_PIPERX4EQDONE (PIPERX4EQDONE_IN, PIPERX4EQDONE);
  buf B_PIPERX4EQLPADAPTDONE (PIPERX4EQLPADAPTDONE_IN, PIPERX4EQLPADAPTDONE);
  buf B_PIPERX4EQLPLFFSSEL (PIPERX4EQLPLFFSSEL_IN, PIPERX4EQLPLFFSSEL);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET0 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[0], PIPERX4EQLPNEWTXCOEFFORPRESET[0]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET1 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[1], PIPERX4EQLPNEWTXCOEFFORPRESET[1]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET10 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[10], PIPERX4EQLPNEWTXCOEFFORPRESET[10]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET11 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[11], PIPERX4EQLPNEWTXCOEFFORPRESET[11]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET12 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[12], PIPERX4EQLPNEWTXCOEFFORPRESET[12]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET13 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[13], PIPERX4EQLPNEWTXCOEFFORPRESET[13]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET14 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[14], PIPERX4EQLPNEWTXCOEFFORPRESET[14]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET15 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[15], PIPERX4EQLPNEWTXCOEFFORPRESET[15]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET16 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[16], PIPERX4EQLPNEWTXCOEFFORPRESET[16]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET17 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[17], PIPERX4EQLPNEWTXCOEFFORPRESET[17]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET2 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[2], PIPERX4EQLPNEWTXCOEFFORPRESET[2]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET3 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[3], PIPERX4EQLPNEWTXCOEFFORPRESET[3]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET4 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[4], PIPERX4EQLPNEWTXCOEFFORPRESET[4]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET5 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[5], PIPERX4EQLPNEWTXCOEFFORPRESET[5]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET6 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[6], PIPERX4EQLPNEWTXCOEFFORPRESET[6]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET7 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[7], PIPERX4EQLPNEWTXCOEFFORPRESET[7]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET8 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[8], PIPERX4EQLPNEWTXCOEFFORPRESET[8]);
  buf B_PIPERX4EQLPNEWTXCOEFFORPRESET9 (PIPERX4EQLPNEWTXCOEFFORPRESET_IN[9], PIPERX4EQLPNEWTXCOEFFORPRESET[9]);
  buf B_PIPERX4PHYSTATUS (PIPERX4PHYSTATUS_IN, PIPERX4PHYSTATUS);
  buf B_PIPERX4STARTBLOCK (PIPERX4STARTBLOCK_IN, PIPERX4STARTBLOCK);
  buf B_PIPERX4STATUS0 (PIPERX4STATUS_IN[0], PIPERX4STATUS[0]);
  buf B_PIPERX4STATUS1 (PIPERX4STATUS_IN[1], PIPERX4STATUS[1]);
  buf B_PIPERX4STATUS2 (PIPERX4STATUS_IN[2], PIPERX4STATUS[2]);
  buf B_PIPERX4SYNCHEADER0 (PIPERX4SYNCHEADER_IN[0], PIPERX4SYNCHEADER[0]);
  buf B_PIPERX4SYNCHEADER1 (PIPERX4SYNCHEADER_IN[1], PIPERX4SYNCHEADER[1]);
  buf B_PIPERX4VALID (PIPERX4VALID_IN, PIPERX4VALID);
  buf B_PIPERX5CHARISK0 (PIPERX5CHARISK_IN[0], PIPERX5CHARISK[0]);
  buf B_PIPERX5CHARISK1 (PIPERX5CHARISK_IN[1], PIPERX5CHARISK[1]);
  buf B_PIPERX5DATA0 (PIPERX5DATA_IN[0], PIPERX5DATA[0]);
  buf B_PIPERX5DATA1 (PIPERX5DATA_IN[1], PIPERX5DATA[1]);
  buf B_PIPERX5DATA10 (PIPERX5DATA_IN[10], PIPERX5DATA[10]);
  buf B_PIPERX5DATA11 (PIPERX5DATA_IN[11], PIPERX5DATA[11]);
  buf B_PIPERX5DATA12 (PIPERX5DATA_IN[12], PIPERX5DATA[12]);
  buf B_PIPERX5DATA13 (PIPERX5DATA_IN[13], PIPERX5DATA[13]);
  buf B_PIPERX5DATA14 (PIPERX5DATA_IN[14], PIPERX5DATA[14]);
  buf B_PIPERX5DATA15 (PIPERX5DATA_IN[15], PIPERX5DATA[15]);
  buf B_PIPERX5DATA16 (PIPERX5DATA_IN[16], PIPERX5DATA[16]);
  buf B_PIPERX5DATA17 (PIPERX5DATA_IN[17], PIPERX5DATA[17]);
  buf B_PIPERX5DATA18 (PIPERX5DATA_IN[18], PIPERX5DATA[18]);
  buf B_PIPERX5DATA19 (PIPERX5DATA_IN[19], PIPERX5DATA[19]);
  buf B_PIPERX5DATA2 (PIPERX5DATA_IN[2], PIPERX5DATA[2]);
  buf B_PIPERX5DATA20 (PIPERX5DATA_IN[20], PIPERX5DATA[20]);
  buf B_PIPERX5DATA21 (PIPERX5DATA_IN[21], PIPERX5DATA[21]);
  buf B_PIPERX5DATA22 (PIPERX5DATA_IN[22], PIPERX5DATA[22]);
  buf B_PIPERX5DATA23 (PIPERX5DATA_IN[23], PIPERX5DATA[23]);
  buf B_PIPERX5DATA24 (PIPERX5DATA_IN[24], PIPERX5DATA[24]);
  buf B_PIPERX5DATA25 (PIPERX5DATA_IN[25], PIPERX5DATA[25]);
  buf B_PIPERX5DATA26 (PIPERX5DATA_IN[26], PIPERX5DATA[26]);
  buf B_PIPERX5DATA27 (PIPERX5DATA_IN[27], PIPERX5DATA[27]);
  buf B_PIPERX5DATA28 (PIPERX5DATA_IN[28], PIPERX5DATA[28]);
  buf B_PIPERX5DATA29 (PIPERX5DATA_IN[29], PIPERX5DATA[29]);
  buf B_PIPERX5DATA3 (PIPERX5DATA_IN[3], PIPERX5DATA[3]);
  buf B_PIPERX5DATA30 (PIPERX5DATA_IN[30], PIPERX5DATA[30]);
  buf B_PIPERX5DATA31 (PIPERX5DATA_IN[31], PIPERX5DATA[31]);
  buf B_PIPERX5DATA4 (PIPERX5DATA_IN[4], PIPERX5DATA[4]);
  buf B_PIPERX5DATA5 (PIPERX5DATA_IN[5], PIPERX5DATA[5]);
  buf B_PIPERX5DATA6 (PIPERX5DATA_IN[6], PIPERX5DATA[6]);
  buf B_PIPERX5DATA7 (PIPERX5DATA_IN[7], PIPERX5DATA[7]);
  buf B_PIPERX5DATA8 (PIPERX5DATA_IN[8], PIPERX5DATA[8]);
  buf B_PIPERX5DATA9 (PIPERX5DATA_IN[9], PIPERX5DATA[9]);
  buf B_PIPERX5DATAVALID (PIPERX5DATAVALID_IN, PIPERX5DATAVALID);
  buf B_PIPERX5ELECIDLE (PIPERX5ELECIDLE_IN, PIPERX5ELECIDLE);
  buf B_PIPERX5EQDONE (PIPERX5EQDONE_IN, PIPERX5EQDONE);
  buf B_PIPERX5EQLPADAPTDONE (PIPERX5EQLPADAPTDONE_IN, PIPERX5EQLPADAPTDONE);
  buf B_PIPERX5EQLPLFFSSEL (PIPERX5EQLPLFFSSEL_IN, PIPERX5EQLPLFFSSEL);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET0 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[0], PIPERX5EQLPNEWTXCOEFFORPRESET[0]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET1 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[1], PIPERX5EQLPNEWTXCOEFFORPRESET[1]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET10 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[10], PIPERX5EQLPNEWTXCOEFFORPRESET[10]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET11 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[11], PIPERX5EQLPNEWTXCOEFFORPRESET[11]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET12 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[12], PIPERX5EQLPNEWTXCOEFFORPRESET[12]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET13 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[13], PIPERX5EQLPNEWTXCOEFFORPRESET[13]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET14 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[14], PIPERX5EQLPNEWTXCOEFFORPRESET[14]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET15 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[15], PIPERX5EQLPNEWTXCOEFFORPRESET[15]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET16 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[16], PIPERX5EQLPNEWTXCOEFFORPRESET[16]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET17 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[17], PIPERX5EQLPNEWTXCOEFFORPRESET[17]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET2 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[2], PIPERX5EQLPNEWTXCOEFFORPRESET[2]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET3 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[3], PIPERX5EQLPNEWTXCOEFFORPRESET[3]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET4 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[4], PIPERX5EQLPNEWTXCOEFFORPRESET[4]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET5 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[5], PIPERX5EQLPNEWTXCOEFFORPRESET[5]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET6 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[6], PIPERX5EQLPNEWTXCOEFFORPRESET[6]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET7 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[7], PIPERX5EQLPNEWTXCOEFFORPRESET[7]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET8 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[8], PIPERX5EQLPNEWTXCOEFFORPRESET[8]);
  buf B_PIPERX5EQLPNEWTXCOEFFORPRESET9 (PIPERX5EQLPNEWTXCOEFFORPRESET_IN[9], PIPERX5EQLPNEWTXCOEFFORPRESET[9]);
  buf B_PIPERX5PHYSTATUS (PIPERX5PHYSTATUS_IN, PIPERX5PHYSTATUS);
  buf B_PIPERX5STARTBLOCK (PIPERX5STARTBLOCK_IN, PIPERX5STARTBLOCK);
  buf B_PIPERX5STATUS0 (PIPERX5STATUS_IN[0], PIPERX5STATUS[0]);
  buf B_PIPERX5STATUS1 (PIPERX5STATUS_IN[1], PIPERX5STATUS[1]);
  buf B_PIPERX5STATUS2 (PIPERX5STATUS_IN[2], PIPERX5STATUS[2]);
  buf B_PIPERX5SYNCHEADER0 (PIPERX5SYNCHEADER_IN[0], PIPERX5SYNCHEADER[0]);
  buf B_PIPERX5SYNCHEADER1 (PIPERX5SYNCHEADER_IN[1], PIPERX5SYNCHEADER[1]);
  buf B_PIPERX5VALID (PIPERX5VALID_IN, PIPERX5VALID);
  buf B_PIPERX6CHARISK0 (PIPERX6CHARISK_IN[0], PIPERX6CHARISK[0]);
  buf B_PIPERX6CHARISK1 (PIPERX6CHARISK_IN[1], PIPERX6CHARISK[1]);
  buf B_PIPERX6DATA0 (PIPERX6DATA_IN[0], PIPERX6DATA[0]);
  buf B_PIPERX6DATA1 (PIPERX6DATA_IN[1], PIPERX6DATA[1]);
  buf B_PIPERX6DATA10 (PIPERX6DATA_IN[10], PIPERX6DATA[10]);
  buf B_PIPERX6DATA11 (PIPERX6DATA_IN[11], PIPERX6DATA[11]);
  buf B_PIPERX6DATA12 (PIPERX6DATA_IN[12], PIPERX6DATA[12]);
  buf B_PIPERX6DATA13 (PIPERX6DATA_IN[13], PIPERX6DATA[13]);
  buf B_PIPERX6DATA14 (PIPERX6DATA_IN[14], PIPERX6DATA[14]);
  buf B_PIPERX6DATA15 (PIPERX6DATA_IN[15], PIPERX6DATA[15]);
  buf B_PIPERX6DATA16 (PIPERX6DATA_IN[16], PIPERX6DATA[16]);
  buf B_PIPERX6DATA17 (PIPERX6DATA_IN[17], PIPERX6DATA[17]);
  buf B_PIPERX6DATA18 (PIPERX6DATA_IN[18], PIPERX6DATA[18]);
  buf B_PIPERX6DATA19 (PIPERX6DATA_IN[19], PIPERX6DATA[19]);
  buf B_PIPERX6DATA2 (PIPERX6DATA_IN[2], PIPERX6DATA[2]);
  buf B_PIPERX6DATA20 (PIPERX6DATA_IN[20], PIPERX6DATA[20]);
  buf B_PIPERX6DATA21 (PIPERX6DATA_IN[21], PIPERX6DATA[21]);
  buf B_PIPERX6DATA22 (PIPERX6DATA_IN[22], PIPERX6DATA[22]);
  buf B_PIPERX6DATA23 (PIPERX6DATA_IN[23], PIPERX6DATA[23]);
  buf B_PIPERX6DATA24 (PIPERX6DATA_IN[24], PIPERX6DATA[24]);
  buf B_PIPERX6DATA25 (PIPERX6DATA_IN[25], PIPERX6DATA[25]);
  buf B_PIPERX6DATA26 (PIPERX6DATA_IN[26], PIPERX6DATA[26]);
  buf B_PIPERX6DATA27 (PIPERX6DATA_IN[27], PIPERX6DATA[27]);
  buf B_PIPERX6DATA28 (PIPERX6DATA_IN[28], PIPERX6DATA[28]);
  buf B_PIPERX6DATA29 (PIPERX6DATA_IN[29], PIPERX6DATA[29]);
  buf B_PIPERX6DATA3 (PIPERX6DATA_IN[3], PIPERX6DATA[3]);
  buf B_PIPERX6DATA30 (PIPERX6DATA_IN[30], PIPERX6DATA[30]);
  buf B_PIPERX6DATA31 (PIPERX6DATA_IN[31], PIPERX6DATA[31]);
  buf B_PIPERX6DATA4 (PIPERX6DATA_IN[4], PIPERX6DATA[4]);
  buf B_PIPERX6DATA5 (PIPERX6DATA_IN[5], PIPERX6DATA[5]);
  buf B_PIPERX6DATA6 (PIPERX6DATA_IN[6], PIPERX6DATA[6]);
  buf B_PIPERX6DATA7 (PIPERX6DATA_IN[7], PIPERX6DATA[7]);
  buf B_PIPERX6DATA8 (PIPERX6DATA_IN[8], PIPERX6DATA[8]);
  buf B_PIPERX6DATA9 (PIPERX6DATA_IN[9], PIPERX6DATA[9]);
  buf B_PIPERX6DATAVALID (PIPERX6DATAVALID_IN, PIPERX6DATAVALID);
  buf B_PIPERX6ELECIDLE (PIPERX6ELECIDLE_IN, PIPERX6ELECIDLE);
  buf B_PIPERX6EQDONE (PIPERX6EQDONE_IN, PIPERX6EQDONE);
  buf B_PIPERX6EQLPADAPTDONE (PIPERX6EQLPADAPTDONE_IN, PIPERX6EQLPADAPTDONE);
  buf B_PIPERX6EQLPLFFSSEL (PIPERX6EQLPLFFSSEL_IN, PIPERX6EQLPLFFSSEL);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET0 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[0], PIPERX6EQLPNEWTXCOEFFORPRESET[0]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET1 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[1], PIPERX6EQLPNEWTXCOEFFORPRESET[1]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET10 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[10], PIPERX6EQLPNEWTXCOEFFORPRESET[10]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET11 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[11], PIPERX6EQLPNEWTXCOEFFORPRESET[11]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET12 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[12], PIPERX6EQLPNEWTXCOEFFORPRESET[12]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET13 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[13], PIPERX6EQLPNEWTXCOEFFORPRESET[13]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET14 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[14], PIPERX6EQLPNEWTXCOEFFORPRESET[14]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET15 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[15], PIPERX6EQLPNEWTXCOEFFORPRESET[15]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET16 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[16], PIPERX6EQLPNEWTXCOEFFORPRESET[16]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET17 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[17], PIPERX6EQLPNEWTXCOEFFORPRESET[17]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET2 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[2], PIPERX6EQLPNEWTXCOEFFORPRESET[2]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET3 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[3], PIPERX6EQLPNEWTXCOEFFORPRESET[3]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET4 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[4], PIPERX6EQLPNEWTXCOEFFORPRESET[4]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET5 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[5], PIPERX6EQLPNEWTXCOEFFORPRESET[5]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET6 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[6], PIPERX6EQLPNEWTXCOEFFORPRESET[6]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET7 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[7], PIPERX6EQLPNEWTXCOEFFORPRESET[7]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET8 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[8], PIPERX6EQLPNEWTXCOEFFORPRESET[8]);
  buf B_PIPERX6EQLPNEWTXCOEFFORPRESET9 (PIPERX6EQLPNEWTXCOEFFORPRESET_IN[9], PIPERX6EQLPNEWTXCOEFFORPRESET[9]);
  buf B_PIPERX6PHYSTATUS (PIPERX6PHYSTATUS_IN, PIPERX6PHYSTATUS);
  buf B_PIPERX6STARTBLOCK (PIPERX6STARTBLOCK_IN, PIPERX6STARTBLOCK);
  buf B_PIPERX6STATUS0 (PIPERX6STATUS_IN[0], PIPERX6STATUS[0]);
  buf B_PIPERX6STATUS1 (PIPERX6STATUS_IN[1], PIPERX6STATUS[1]);
  buf B_PIPERX6STATUS2 (PIPERX6STATUS_IN[2], PIPERX6STATUS[2]);
  buf B_PIPERX6SYNCHEADER0 (PIPERX6SYNCHEADER_IN[0], PIPERX6SYNCHEADER[0]);
  buf B_PIPERX6SYNCHEADER1 (PIPERX6SYNCHEADER_IN[1], PIPERX6SYNCHEADER[1]);
  buf B_PIPERX6VALID (PIPERX6VALID_IN, PIPERX6VALID);
  buf B_PIPERX7CHARISK0 (PIPERX7CHARISK_IN[0], PIPERX7CHARISK[0]);
  buf B_PIPERX7CHARISK1 (PIPERX7CHARISK_IN[1], PIPERX7CHARISK[1]);
  buf B_PIPERX7DATA0 (PIPERX7DATA_IN[0], PIPERX7DATA[0]);
  buf B_PIPERX7DATA1 (PIPERX7DATA_IN[1], PIPERX7DATA[1]);
  buf B_PIPERX7DATA10 (PIPERX7DATA_IN[10], PIPERX7DATA[10]);
  buf B_PIPERX7DATA11 (PIPERX7DATA_IN[11], PIPERX7DATA[11]);
  buf B_PIPERX7DATA12 (PIPERX7DATA_IN[12], PIPERX7DATA[12]);
  buf B_PIPERX7DATA13 (PIPERX7DATA_IN[13], PIPERX7DATA[13]);
  buf B_PIPERX7DATA14 (PIPERX7DATA_IN[14], PIPERX7DATA[14]);
  buf B_PIPERX7DATA15 (PIPERX7DATA_IN[15], PIPERX7DATA[15]);
  buf B_PIPERX7DATA16 (PIPERX7DATA_IN[16], PIPERX7DATA[16]);
  buf B_PIPERX7DATA17 (PIPERX7DATA_IN[17], PIPERX7DATA[17]);
  buf B_PIPERX7DATA18 (PIPERX7DATA_IN[18], PIPERX7DATA[18]);
  buf B_PIPERX7DATA19 (PIPERX7DATA_IN[19], PIPERX7DATA[19]);
  buf B_PIPERX7DATA2 (PIPERX7DATA_IN[2], PIPERX7DATA[2]);
  buf B_PIPERX7DATA20 (PIPERX7DATA_IN[20], PIPERX7DATA[20]);
  buf B_PIPERX7DATA21 (PIPERX7DATA_IN[21], PIPERX7DATA[21]);
  buf B_PIPERX7DATA22 (PIPERX7DATA_IN[22], PIPERX7DATA[22]);
  buf B_PIPERX7DATA23 (PIPERX7DATA_IN[23], PIPERX7DATA[23]);
  buf B_PIPERX7DATA24 (PIPERX7DATA_IN[24], PIPERX7DATA[24]);
  buf B_PIPERX7DATA25 (PIPERX7DATA_IN[25], PIPERX7DATA[25]);
  buf B_PIPERX7DATA26 (PIPERX7DATA_IN[26], PIPERX7DATA[26]);
  buf B_PIPERX7DATA27 (PIPERX7DATA_IN[27], PIPERX7DATA[27]);
  buf B_PIPERX7DATA28 (PIPERX7DATA_IN[28], PIPERX7DATA[28]);
  buf B_PIPERX7DATA29 (PIPERX7DATA_IN[29], PIPERX7DATA[29]);
  buf B_PIPERX7DATA3 (PIPERX7DATA_IN[3], PIPERX7DATA[3]);
  buf B_PIPERX7DATA30 (PIPERX7DATA_IN[30], PIPERX7DATA[30]);
  buf B_PIPERX7DATA31 (PIPERX7DATA_IN[31], PIPERX7DATA[31]);
  buf B_PIPERX7DATA4 (PIPERX7DATA_IN[4], PIPERX7DATA[4]);
  buf B_PIPERX7DATA5 (PIPERX7DATA_IN[5], PIPERX7DATA[5]);
  buf B_PIPERX7DATA6 (PIPERX7DATA_IN[6], PIPERX7DATA[6]);
  buf B_PIPERX7DATA7 (PIPERX7DATA_IN[7], PIPERX7DATA[7]);
  buf B_PIPERX7DATA8 (PIPERX7DATA_IN[8], PIPERX7DATA[8]);
  buf B_PIPERX7DATA9 (PIPERX7DATA_IN[9], PIPERX7DATA[9]);
  buf B_PIPERX7DATAVALID (PIPERX7DATAVALID_IN, PIPERX7DATAVALID);
  buf B_PIPERX7ELECIDLE (PIPERX7ELECIDLE_IN, PIPERX7ELECIDLE);
  buf B_PIPERX7EQDONE (PIPERX7EQDONE_IN, PIPERX7EQDONE);
  buf B_PIPERX7EQLPADAPTDONE (PIPERX7EQLPADAPTDONE_IN, PIPERX7EQLPADAPTDONE);
  buf B_PIPERX7EQLPLFFSSEL (PIPERX7EQLPLFFSSEL_IN, PIPERX7EQLPLFFSSEL);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET0 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[0], PIPERX7EQLPNEWTXCOEFFORPRESET[0]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET1 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[1], PIPERX7EQLPNEWTXCOEFFORPRESET[1]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET10 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[10], PIPERX7EQLPNEWTXCOEFFORPRESET[10]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET11 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[11], PIPERX7EQLPNEWTXCOEFFORPRESET[11]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET12 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[12], PIPERX7EQLPNEWTXCOEFFORPRESET[12]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET13 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[13], PIPERX7EQLPNEWTXCOEFFORPRESET[13]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET14 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[14], PIPERX7EQLPNEWTXCOEFFORPRESET[14]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET15 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[15], PIPERX7EQLPNEWTXCOEFFORPRESET[15]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET16 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[16], PIPERX7EQLPNEWTXCOEFFORPRESET[16]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET17 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[17], PIPERX7EQLPNEWTXCOEFFORPRESET[17]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET2 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[2], PIPERX7EQLPNEWTXCOEFFORPRESET[2]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET3 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[3], PIPERX7EQLPNEWTXCOEFFORPRESET[3]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET4 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[4], PIPERX7EQLPNEWTXCOEFFORPRESET[4]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET5 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[5], PIPERX7EQLPNEWTXCOEFFORPRESET[5]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET6 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[6], PIPERX7EQLPNEWTXCOEFFORPRESET[6]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET7 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[7], PIPERX7EQLPNEWTXCOEFFORPRESET[7]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET8 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[8], PIPERX7EQLPNEWTXCOEFFORPRESET[8]);
  buf B_PIPERX7EQLPNEWTXCOEFFORPRESET9 (PIPERX7EQLPNEWTXCOEFFORPRESET_IN[9], PIPERX7EQLPNEWTXCOEFFORPRESET[9]);
  buf B_PIPERX7PHYSTATUS (PIPERX7PHYSTATUS_IN, PIPERX7PHYSTATUS);
  buf B_PIPERX7STARTBLOCK (PIPERX7STARTBLOCK_IN, PIPERX7STARTBLOCK);
  buf B_PIPERX7STATUS0 (PIPERX7STATUS_IN[0], PIPERX7STATUS[0]);
  buf B_PIPERX7STATUS1 (PIPERX7STATUS_IN[1], PIPERX7STATUS[1]);
  buf B_PIPERX7STATUS2 (PIPERX7STATUS_IN[2], PIPERX7STATUS[2]);
  buf B_PIPERX7SYNCHEADER0 (PIPERX7SYNCHEADER_IN[0], PIPERX7SYNCHEADER[0]);
  buf B_PIPERX7SYNCHEADER1 (PIPERX7SYNCHEADER_IN[1], PIPERX7SYNCHEADER[1]);
  buf B_PIPERX7VALID (PIPERX7VALID_IN, PIPERX7VALID);
  buf B_PIPETX0EQCOEFF0 (PIPETX0EQCOEFF_IN[0], PIPETX0EQCOEFF[0]);
  buf B_PIPETX0EQCOEFF1 (PIPETX0EQCOEFF_IN[1], PIPETX0EQCOEFF[1]);
  buf B_PIPETX0EQCOEFF10 (PIPETX0EQCOEFF_IN[10], PIPETX0EQCOEFF[10]);
  buf B_PIPETX0EQCOEFF11 (PIPETX0EQCOEFF_IN[11], PIPETX0EQCOEFF[11]);
  buf B_PIPETX0EQCOEFF12 (PIPETX0EQCOEFF_IN[12], PIPETX0EQCOEFF[12]);
  buf B_PIPETX0EQCOEFF13 (PIPETX0EQCOEFF_IN[13], PIPETX0EQCOEFF[13]);
  buf B_PIPETX0EQCOEFF14 (PIPETX0EQCOEFF_IN[14], PIPETX0EQCOEFF[14]);
  buf B_PIPETX0EQCOEFF15 (PIPETX0EQCOEFF_IN[15], PIPETX0EQCOEFF[15]);
  buf B_PIPETX0EQCOEFF16 (PIPETX0EQCOEFF_IN[16], PIPETX0EQCOEFF[16]);
  buf B_PIPETX0EQCOEFF17 (PIPETX0EQCOEFF_IN[17], PIPETX0EQCOEFF[17]);
  buf B_PIPETX0EQCOEFF2 (PIPETX0EQCOEFF_IN[2], PIPETX0EQCOEFF[2]);
  buf B_PIPETX0EQCOEFF3 (PIPETX0EQCOEFF_IN[3], PIPETX0EQCOEFF[3]);
  buf B_PIPETX0EQCOEFF4 (PIPETX0EQCOEFF_IN[4], PIPETX0EQCOEFF[4]);
  buf B_PIPETX0EQCOEFF5 (PIPETX0EQCOEFF_IN[5], PIPETX0EQCOEFF[5]);
  buf B_PIPETX0EQCOEFF6 (PIPETX0EQCOEFF_IN[6], PIPETX0EQCOEFF[6]);
  buf B_PIPETX0EQCOEFF7 (PIPETX0EQCOEFF_IN[7], PIPETX0EQCOEFF[7]);
  buf B_PIPETX0EQCOEFF8 (PIPETX0EQCOEFF_IN[8], PIPETX0EQCOEFF[8]);
  buf B_PIPETX0EQCOEFF9 (PIPETX0EQCOEFF_IN[9], PIPETX0EQCOEFF[9]);
  buf B_PIPETX0EQDONE (PIPETX0EQDONE_IN, PIPETX0EQDONE);
  buf B_PIPETX1EQCOEFF0 (PIPETX1EQCOEFF_IN[0], PIPETX1EQCOEFF[0]);
  buf B_PIPETX1EQCOEFF1 (PIPETX1EQCOEFF_IN[1], PIPETX1EQCOEFF[1]);
  buf B_PIPETX1EQCOEFF10 (PIPETX1EQCOEFF_IN[10], PIPETX1EQCOEFF[10]);
  buf B_PIPETX1EQCOEFF11 (PIPETX1EQCOEFF_IN[11], PIPETX1EQCOEFF[11]);
  buf B_PIPETX1EQCOEFF12 (PIPETX1EQCOEFF_IN[12], PIPETX1EQCOEFF[12]);
  buf B_PIPETX1EQCOEFF13 (PIPETX1EQCOEFF_IN[13], PIPETX1EQCOEFF[13]);
  buf B_PIPETX1EQCOEFF14 (PIPETX1EQCOEFF_IN[14], PIPETX1EQCOEFF[14]);
  buf B_PIPETX1EQCOEFF15 (PIPETX1EQCOEFF_IN[15], PIPETX1EQCOEFF[15]);
  buf B_PIPETX1EQCOEFF16 (PIPETX1EQCOEFF_IN[16], PIPETX1EQCOEFF[16]);
  buf B_PIPETX1EQCOEFF17 (PIPETX1EQCOEFF_IN[17], PIPETX1EQCOEFF[17]);
  buf B_PIPETX1EQCOEFF2 (PIPETX1EQCOEFF_IN[2], PIPETX1EQCOEFF[2]);
  buf B_PIPETX1EQCOEFF3 (PIPETX1EQCOEFF_IN[3], PIPETX1EQCOEFF[3]);
  buf B_PIPETX1EQCOEFF4 (PIPETX1EQCOEFF_IN[4], PIPETX1EQCOEFF[4]);
  buf B_PIPETX1EQCOEFF5 (PIPETX1EQCOEFF_IN[5], PIPETX1EQCOEFF[5]);
  buf B_PIPETX1EQCOEFF6 (PIPETX1EQCOEFF_IN[6], PIPETX1EQCOEFF[6]);
  buf B_PIPETX1EQCOEFF7 (PIPETX1EQCOEFF_IN[7], PIPETX1EQCOEFF[7]);
  buf B_PIPETX1EQCOEFF8 (PIPETX1EQCOEFF_IN[8], PIPETX1EQCOEFF[8]);
  buf B_PIPETX1EQCOEFF9 (PIPETX1EQCOEFF_IN[9], PIPETX1EQCOEFF[9]);
  buf B_PIPETX1EQDONE (PIPETX1EQDONE_IN, PIPETX1EQDONE);
  buf B_PIPETX2EQCOEFF0 (PIPETX2EQCOEFF_IN[0], PIPETX2EQCOEFF[0]);
  buf B_PIPETX2EQCOEFF1 (PIPETX2EQCOEFF_IN[1], PIPETX2EQCOEFF[1]);
  buf B_PIPETX2EQCOEFF10 (PIPETX2EQCOEFF_IN[10], PIPETX2EQCOEFF[10]);
  buf B_PIPETX2EQCOEFF11 (PIPETX2EQCOEFF_IN[11], PIPETX2EQCOEFF[11]);
  buf B_PIPETX2EQCOEFF12 (PIPETX2EQCOEFF_IN[12], PIPETX2EQCOEFF[12]);
  buf B_PIPETX2EQCOEFF13 (PIPETX2EQCOEFF_IN[13], PIPETX2EQCOEFF[13]);
  buf B_PIPETX2EQCOEFF14 (PIPETX2EQCOEFF_IN[14], PIPETX2EQCOEFF[14]);
  buf B_PIPETX2EQCOEFF15 (PIPETX2EQCOEFF_IN[15], PIPETX2EQCOEFF[15]);
  buf B_PIPETX2EQCOEFF16 (PIPETX2EQCOEFF_IN[16], PIPETX2EQCOEFF[16]);
  buf B_PIPETX2EQCOEFF17 (PIPETX2EQCOEFF_IN[17], PIPETX2EQCOEFF[17]);
  buf B_PIPETX2EQCOEFF2 (PIPETX2EQCOEFF_IN[2], PIPETX2EQCOEFF[2]);
  buf B_PIPETX2EQCOEFF3 (PIPETX2EQCOEFF_IN[3], PIPETX2EQCOEFF[3]);
  buf B_PIPETX2EQCOEFF4 (PIPETX2EQCOEFF_IN[4], PIPETX2EQCOEFF[4]);
  buf B_PIPETX2EQCOEFF5 (PIPETX2EQCOEFF_IN[5], PIPETX2EQCOEFF[5]);
  buf B_PIPETX2EQCOEFF6 (PIPETX2EQCOEFF_IN[6], PIPETX2EQCOEFF[6]);
  buf B_PIPETX2EQCOEFF7 (PIPETX2EQCOEFF_IN[7], PIPETX2EQCOEFF[7]);
  buf B_PIPETX2EQCOEFF8 (PIPETX2EQCOEFF_IN[8], PIPETX2EQCOEFF[8]);
  buf B_PIPETX2EQCOEFF9 (PIPETX2EQCOEFF_IN[9], PIPETX2EQCOEFF[9]);
  buf B_PIPETX2EQDONE (PIPETX2EQDONE_IN, PIPETX2EQDONE);
  buf B_PIPETX3EQCOEFF0 (PIPETX3EQCOEFF_IN[0], PIPETX3EQCOEFF[0]);
  buf B_PIPETX3EQCOEFF1 (PIPETX3EQCOEFF_IN[1], PIPETX3EQCOEFF[1]);
  buf B_PIPETX3EQCOEFF10 (PIPETX3EQCOEFF_IN[10], PIPETX3EQCOEFF[10]);
  buf B_PIPETX3EQCOEFF11 (PIPETX3EQCOEFF_IN[11], PIPETX3EQCOEFF[11]);
  buf B_PIPETX3EQCOEFF12 (PIPETX3EQCOEFF_IN[12], PIPETX3EQCOEFF[12]);
  buf B_PIPETX3EQCOEFF13 (PIPETX3EQCOEFF_IN[13], PIPETX3EQCOEFF[13]);
  buf B_PIPETX3EQCOEFF14 (PIPETX3EQCOEFF_IN[14], PIPETX3EQCOEFF[14]);
  buf B_PIPETX3EQCOEFF15 (PIPETX3EQCOEFF_IN[15], PIPETX3EQCOEFF[15]);
  buf B_PIPETX3EQCOEFF16 (PIPETX3EQCOEFF_IN[16], PIPETX3EQCOEFF[16]);
  buf B_PIPETX3EQCOEFF17 (PIPETX3EQCOEFF_IN[17], PIPETX3EQCOEFF[17]);
  buf B_PIPETX3EQCOEFF2 (PIPETX3EQCOEFF_IN[2], PIPETX3EQCOEFF[2]);
  buf B_PIPETX3EQCOEFF3 (PIPETX3EQCOEFF_IN[3], PIPETX3EQCOEFF[3]);
  buf B_PIPETX3EQCOEFF4 (PIPETX3EQCOEFF_IN[4], PIPETX3EQCOEFF[4]);
  buf B_PIPETX3EQCOEFF5 (PIPETX3EQCOEFF_IN[5], PIPETX3EQCOEFF[5]);
  buf B_PIPETX3EQCOEFF6 (PIPETX3EQCOEFF_IN[6], PIPETX3EQCOEFF[6]);
  buf B_PIPETX3EQCOEFF7 (PIPETX3EQCOEFF_IN[7], PIPETX3EQCOEFF[7]);
  buf B_PIPETX3EQCOEFF8 (PIPETX3EQCOEFF_IN[8], PIPETX3EQCOEFF[8]);
  buf B_PIPETX3EQCOEFF9 (PIPETX3EQCOEFF_IN[9], PIPETX3EQCOEFF[9]);
  buf B_PIPETX3EQDONE (PIPETX3EQDONE_IN, PIPETX3EQDONE);
  buf B_PIPETX4EQCOEFF0 (PIPETX4EQCOEFF_IN[0], PIPETX4EQCOEFF[0]);
  buf B_PIPETX4EQCOEFF1 (PIPETX4EQCOEFF_IN[1], PIPETX4EQCOEFF[1]);
  buf B_PIPETX4EQCOEFF10 (PIPETX4EQCOEFF_IN[10], PIPETX4EQCOEFF[10]);
  buf B_PIPETX4EQCOEFF11 (PIPETX4EQCOEFF_IN[11], PIPETX4EQCOEFF[11]);
  buf B_PIPETX4EQCOEFF12 (PIPETX4EQCOEFF_IN[12], PIPETX4EQCOEFF[12]);
  buf B_PIPETX4EQCOEFF13 (PIPETX4EQCOEFF_IN[13], PIPETX4EQCOEFF[13]);
  buf B_PIPETX4EQCOEFF14 (PIPETX4EQCOEFF_IN[14], PIPETX4EQCOEFF[14]);
  buf B_PIPETX4EQCOEFF15 (PIPETX4EQCOEFF_IN[15], PIPETX4EQCOEFF[15]);
  buf B_PIPETX4EQCOEFF16 (PIPETX4EQCOEFF_IN[16], PIPETX4EQCOEFF[16]);
  buf B_PIPETX4EQCOEFF17 (PIPETX4EQCOEFF_IN[17], PIPETX4EQCOEFF[17]);
  buf B_PIPETX4EQCOEFF2 (PIPETX4EQCOEFF_IN[2], PIPETX4EQCOEFF[2]);
  buf B_PIPETX4EQCOEFF3 (PIPETX4EQCOEFF_IN[3], PIPETX4EQCOEFF[3]);
  buf B_PIPETX4EQCOEFF4 (PIPETX4EQCOEFF_IN[4], PIPETX4EQCOEFF[4]);
  buf B_PIPETX4EQCOEFF5 (PIPETX4EQCOEFF_IN[5], PIPETX4EQCOEFF[5]);
  buf B_PIPETX4EQCOEFF6 (PIPETX4EQCOEFF_IN[6], PIPETX4EQCOEFF[6]);
  buf B_PIPETX4EQCOEFF7 (PIPETX4EQCOEFF_IN[7], PIPETX4EQCOEFF[7]);
  buf B_PIPETX4EQCOEFF8 (PIPETX4EQCOEFF_IN[8], PIPETX4EQCOEFF[8]);
  buf B_PIPETX4EQCOEFF9 (PIPETX4EQCOEFF_IN[9], PIPETX4EQCOEFF[9]);
  buf B_PIPETX4EQDONE (PIPETX4EQDONE_IN, PIPETX4EQDONE);
  buf B_PIPETX5EQCOEFF0 (PIPETX5EQCOEFF_IN[0], PIPETX5EQCOEFF[0]);
  buf B_PIPETX5EQCOEFF1 (PIPETX5EQCOEFF_IN[1], PIPETX5EQCOEFF[1]);
  buf B_PIPETX5EQCOEFF10 (PIPETX5EQCOEFF_IN[10], PIPETX5EQCOEFF[10]);
  buf B_PIPETX5EQCOEFF11 (PIPETX5EQCOEFF_IN[11], PIPETX5EQCOEFF[11]);
  buf B_PIPETX5EQCOEFF12 (PIPETX5EQCOEFF_IN[12], PIPETX5EQCOEFF[12]);
  buf B_PIPETX5EQCOEFF13 (PIPETX5EQCOEFF_IN[13], PIPETX5EQCOEFF[13]);
  buf B_PIPETX5EQCOEFF14 (PIPETX5EQCOEFF_IN[14], PIPETX5EQCOEFF[14]);
  buf B_PIPETX5EQCOEFF15 (PIPETX5EQCOEFF_IN[15], PIPETX5EQCOEFF[15]);
  buf B_PIPETX5EQCOEFF16 (PIPETX5EQCOEFF_IN[16], PIPETX5EQCOEFF[16]);
  buf B_PIPETX5EQCOEFF17 (PIPETX5EQCOEFF_IN[17], PIPETX5EQCOEFF[17]);
  buf B_PIPETX5EQCOEFF2 (PIPETX5EQCOEFF_IN[2], PIPETX5EQCOEFF[2]);
  buf B_PIPETX5EQCOEFF3 (PIPETX5EQCOEFF_IN[3], PIPETX5EQCOEFF[3]);
  buf B_PIPETX5EQCOEFF4 (PIPETX5EQCOEFF_IN[4], PIPETX5EQCOEFF[4]);
  buf B_PIPETX5EQCOEFF5 (PIPETX5EQCOEFF_IN[5], PIPETX5EQCOEFF[5]);
  buf B_PIPETX5EQCOEFF6 (PIPETX5EQCOEFF_IN[6], PIPETX5EQCOEFF[6]);
  buf B_PIPETX5EQCOEFF7 (PIPETX5EQCOEFF_IN[7], PIPETX5EQCOEFF[7]);
  buf B_PIPETX5EQCOEFF8 (PIPETX5EQCOEFF_IN[8], PIPETX5EQCOEFF[8]);
  buf B_PIPETX5EQCOEFF9 (PIPETX5EQCOEFF_IN[9], PIPETX5EQCOEFF[9]);
  buf B_PIPETX5EQDONE (PIPETX5EQDONE_IN, PIPETX5EQDONE);
  buf B_PIPETX6EQCOEFF0 (PIPETX6EQCOEFF_IN[0], PIPETX6EQCOEFF[0]);
  buf B_PIPETX6EQCOEFF1 (PIPETX6EQCOEFF_IN[1], PIPETX6EQCOEFF[1]);
  buf B_PIPETX6EQCOEFF10 (PIPETX6EQCOEFF_IN[10], PIPETX6EQCOEFF[10]);
  buf B_PIPETX6EQCOEFF11 (PIPETX6EQCOEFF_IN[11], PIPETX6EQCOEFF[11]);
  buf B_PIPETX6EQCOEFF12 (PIPETX6EQCOEFF_IN[12], PIPETX6EQCOEFF[12]);
  buf B_PIPETX6EQCOEFF13 (PIPETX6EQCOEFF_IN[13], PIPETX6EQCOEFF[13]);
  buf B_PIPETX6EQCOEFF14 (PIPETX6EQCOEFF_IN[14], PIPETX6EQCOEFF[14]);
  buf B_PIPETX6EQCOEFF15 (PIPETX6EQCOEFF_IN[15], PIPETX6EQCOEFF[15]);
  buf B_PIPETX6EQCOEFF16 (PIPETX6EQCOEFF_IN[16], PIPETX6EQCOEFF[16]);
  buf B_PIPETX6EQCOEFF17 (PIPETX6EQCOEFF_IN[17], PIPETX6EQCOEFF[17]);
  buf B_PIPETX6EQCOEFF2 (PIPETX6EQCOEFF_IN[2], PIPETX6EQCOEFF[2]);
  buf B_PIPETX6EQCOEFF3 (PIPETX6EQCOEFF_IN[3], PIPETX6EQCOEFF[3]);
  buf B_PIPETX6EQCOEFF4 (PIPETX6EQCOEFF_IN[4], PIPETX6EQCOEFF[4]);
  buf B_PIPETX6EQCOEFF5 (PIPETX6EQCOEFF_IN[5], PIPETX6EQCOEFF[5]);
  buf B_PIPETX6EQCOEFF6 (PIPETX6EQCOEFF_IN[6], PIPETX6EQCOEFF[6]);
  buf B_PIPETX6EQCOEFF7 (PIPETX6EQCOEFF_IN[7], PIPETX6EQCOEFF[7]);
  buf B_PIPETX6EQCOEFF8 (PIPETX6EQCOEFF_IN[8], PIPETX6EQCOEFF[8]);
  buf B_PIPETX6EQCOEFF9 (PIPETX6EQCOEFF_IN[9], PIPETX6EQCOEFF[9]);
  buf B_PIPETX6EQDONE (PIPETX6EQDONE_IN, PIPETX6EQDONE);
  buf B_PIPETX7EQCOEFF0 (PIPETX7EQCOEFF_IN[0], PIPETX7EQCOEFF[0]);
  buf B_PIPETX7EQCOEFF1 (PIPETX7EQCOEFF_IN[1], PIPETX7EQCOEFF[1]);
  buf B_PIPETX7EQCOEFF10 (PIPETX7EQCOEFF_IN[10], PIPETX7EQCOEFF[10]);
  buf B_PIPETX7EQCOEFF11 (PIPETX7EQCOEFF_IN[11], PIPETX7EQCOEFF[11]);
  buf B_PIPETX7EQCOEFF12 (PIPETX7EQCOEFF_IN[12], PIPETX7EQCOEFF[12]);
  buf B_PIPETX7EQCOEFF13 (PIPETX7EQCOEFF_IN[13], PIPETX7EQCOEFF[13]);
  buf B_PIPETX7EQCOEFF14 (PIPETX7EQCOEFF_IN[14], PIPETX7EQCOEFF[14]);
  buf B_PIPETX7EQCOEFF15 (PIPETX7EQCOEFF_IN[15], PIPETX7EQCOEFF[15]);
  buf B_PIPETX7EQCOEFF16 (PIPETX7EQCOEFF_IN[16], PIPETX7EQCOEFF[16]);
  buf B_PIPETX7EQCOEFF17 (PIPETX7EQCOEFF_IN[17], PIPETX7EQCOEFF[17]);
  buf B_PIPETX7EQCOEFF2 (PIPETX7EQCOEFF_IN[2], PIPETX7EQCOEFF[2]);
  buf B_PIPETX7EQCOEFF3 (PIPETX7EQCOEFF_IN[3], PIPETX7EQCOEFF[3]);
  buf B_PIPETX7EQCOEFF4 (PIPETX7EQCOEFF_IN[4], PIPETX7EQCOEFF[4]);
  buf B_PIPETX7EQCOEFF5 (PIPETX7EQCOEFF_IN[5], PIPETX7EQCOEFF[5]);
  buf B_PIPETX7EQCOEFF6 (PIPETX7EQCOEFF_IN[6], PIPETX7EQCOEFF[6]);
  buf B_PIPETX7EQCOEFF7 (PIPETX7EQCOEFF_IN[7], PIPETX7EQCOEFF[7]);
  buf B_PIPETX7EQCOEFF8 (PIPETX7EQCOEFF_IN[8], PIPETX7EQCOEFF[8]);
  buf B_PIPETX7EQCOEFF9 (PIPETX7EQCOEFF_IN[9], PIPETX7EQCOEFF[9]);
  buf B_PIPETX7EQDONE (PIPETX7EQDONE_IN, PIPETX7EQDONE);
  buf B_PLDISABLESCRAMBLER (PLDISABLESCRAMBLER_IN, PLDISABLESCRAMBLER);
  buf B_PLEQRESETEIEOSCOUNT (PLEQRESETEIEOSCOUNT_IN, PLEQRESETEIEOSCOUNT);
  buf B_PLGEN3PCSDISABLE (PLGEN3PCSDISABLE_IN, PLGEN3PCSDISABLE);
  buf B_PLGEN3PCSRXSYNCDONE0 (PLGEN3PCSRXSYNCDONE_IN[0], PLGEN3PCSRXSYNCDONE[0]);
  buf B_PLGEN3PCSRXSYNCDONE1 (PLGEN3PCSRXSYNCDONE_IN[1], PLGEN3PCSRXSYNCDONE[1]);
  buf B_PLGEN3PCSRXSYNCDONE2 (PLGEN3PCSRXSYNCDONE_IN[2], PLGEN3PCSRXSYNCDONE[2]);
  buf B_PLGEN3PCSRXSYNCDONE3 (PLGEN3PCSRXSYNCDONE_IN[3], PLGEN3PCSRXSYNCDONE[3]);
  buf B_PLGEN3PCSRXSYNCDONE4 (PLGEN3PCSRXSYNCDONE_IN[4], PLGEN3PCSRXSYNCDONE[4]);
  buf B_PLGEN3PCSRXSYNCDONE5 (PLGEN3PCSRXSYNCDONE_IN[5], PLGEN3PCSRXSYNCDONE[5]);
  buf B_PLGEN3PCSRXSYNCDONE6 (PLGEN3PCSRXSYNCDONE_IN[6], PLGEN3PCSRXSYNCDONE[6]);
  buf B_PLGEN3PCSRXSYNCDONE7 (PLGEN3PCSRXSYNCDONE_IN[7], PLGEN3PCSRXSYNCDONE[7]);
  buf B_RECCLK (RECCLK_IN, RECCLK);
  buf B_RESETN (RESETN_IN, RESETN);
  buf B_SAXISCCTDATA0 (SAXISCCTDATA_IN[0], SAXISCCTDATA[0]);
  buf B_SAXISCCTDATA1 (SAXISCCTDATA_IN[1], SAXISCCTDATA[1]);
  buf B_SAXISCCTDATA10 (SAXISCCTDATA_IN[10], SAXISCCTDATA[10]);
  buf B_SAXISCCTDATA100 (SAXISCCTDATA_IN[100], SAXISCCTDATA[100]);
  buf B_SAXISCCTDATA101 (SAXISCCTDATA_IN[101], SAXISCCTDATA[101]);
  buf B_SAXISCCTDATA102 (SAXISCCTDATA_IN[102], SAXISCCTDATA[102]);
  buf B_SAXISCCTDATA103 (SAXISCCTDATA_IN[103], SAXISCCTDATA[103]);
  buf B_SAXISCCTDATA104 (SAXISCCTDATA_IN[104], SAXISCCTDATA[104]);
  buf B_SAXISCCTDATA105 (SAXISCCTDATA_IN[105], SAXISCCTDATA[105]);
  buf B_SAXISCCTDATA106 (SAXISCCTDATA_IN[106], SAXISCCTDATA[106]);
  buf B_SAXISCCTDATA107 (SAXISCCTDATA_IN[107], SAXISCCTDATA[107]);
  buf B_SAXISCCTDATA108 (SAXISCCTDATA_IN[108], SAXISCCTDATA[108]);
  buf B_SAXISCCTDATA109 (SAXISCCTDATA_IN[109], SAXISCCTDATA[109]);
  buf B_SAXISCCTDATA11 (SAXISCCTDATA_IN[11], SAXISCCTDATA[11]);
  buf B_SAXISCCTDATA110 (SAXISCCTDATA_IN[110], SAXISCCTDATA[110]);
  buf B_SAXISCCTDATA111 (SAXISCCTDATA_IN[111], SAXISCCTDATA[111]);
  buf B_SAXISCCTDATA112 (SAXISCCTDATA_IN[112], SAXISCCTDATA[112]);
  buf B_SAXISCCTDATA113 (SAXISCCTDATA_IN[113], SAXISCCTDATA[113]);
  buf B_SAXISCCTDATA114 (SAXISCCTDATA_IN[114], SAXISCCTDATA[114]);
  buf B_SAXISCCTDATA115 (SAXISCCTDATA_IN[115], SAXISCCTDATA[115]);
  buf B_SAXISCCTDATA116 (SAXISCCTDATA_IN[116], SAXISCCTDATA[116]);
  buf B_SAXISCCTDATA117 (SAXISCCTDATA_IN[117], SAXISCCTDATA[117]);
  buf B_SAXISCCTDATA118 (SAXISCCTDATA_IN[118], SAXISCCTDATA[118]);
  buf B_SAXISCCTDATA119 (SAXISCCTDATA_IN[119], SAXISCCTDATA[119]);
  buf B_SAXISCCTDATA12 (SAXISCCTDATA_IN[12], SAXISCCTDATA[12]);
  buf B_SAXISCCTDATA120 (SAXISCCTDATA_IN[120], SAXISCCTDATA[120]);
  buf B_SAXISCCTDATA121 (SAXISCCTDATA_IN[121], SAXISCCTDATA[121]);
  buf B_SAXISCCTDATA122 (SAXISCCTDATA_IN[122], SAXISCCTDATA[122]);
  buf B_SAXISCCTDATA123 (SAXISCCTDATA_IN[123], SAXISCCTDATA[123]);
  buf B_SAXISCCTDATA124 (SAXISCCTDATA_IN[124], SAXISCCTDATA[124]);
  buf B_SAXISCCTDATA125 (SAXISCCTDATA_IN[125], SAXISCCTDATA[125]);
  buf B_SAXISCCTDATA126 (SAXISCCTDATA_IN[126], SAXISCCTDATA[126]);
  buf B_SAXISCCTDATA127 (SAXISCCTDATA_IN[127], SAXISCCTDATA[127]);
  buf B_SAXISCCTDATA128 (SAXISCCTDATA_IN[128], SAXISCCTDATA[128]);
  buf B_SAXISCCTDATA129 (SAXISCCTDATA_IN[129], SAXISCCTDATA[129]);
  buf B_SAXISCCTDATA13 (SAXISCCTDATA_IN[13], SAXISCCTDATA[13]);
  buf B_SAXISCCTDATA130 (SAXISCCTDATA_IN[130], SAXISCCTDATA[130]);
  buf B_SAXISCCTDATA131 (SAXISCCTDATA_IN[131], SAXISCCTDATA[131]);
  buf B_SAXISCCTDATA132 (SAXISCCTDATA_IN[132], SAXISCCTDATA[132]);
  buf B_SAXISCCTDATA133 (SAXISCCTDATA_IN[133], SAXISCCTDATA[133]);
  buf B_SAXISCCTDATA134 (SAXISCCTDATA_IN[134], SAXISCCTDATA[134]);
  buf B_SAXISCCTDATA135 (SAXISCCTDATA_IN[135], SAXISCCTDATA[135]);
  buf B_SAXISCCTDATA136 (SAXISCCTDATA_IN[136], SAXISCCTDATA[136]);
  buf B_SAXISCCTDATA137 (SAXISCCTDATA_IN[137], SAXISCCTDATA[137]);
  buf B_SAXISCCTDATA138 (SAXISCCTDATA_IN[138], SAXISCCTDATA[138]);
  buf B_SAXISCCTDATA139 (SAXISCCTDATA_IN[139], SAXISCCTDATA[139]);
  buf B_SAXISCCTDATA14 (SAXISCCTDATA_IN[14], SAXISCCTDATA[14]);
  buf B_SAXISCCTDATA140 (SAXISCCTDATA_IN[140], SAXISCCTDATA[140]);
  buf B_SAXISCCTDATA141 (SAXISCCTDATA_IN[141], SAXISCCTDATA[141]);
  buf B_SAXISCCTDATA142 (SAXISCCTDATA_IN[142], SAXISCCTDATA[142]);
  buf B_SAXISCCTDATA143 (SAXISCCTDATA_IN[143], SAXISCCTDATA[143]);
  buf B_SAXISCCTDATA144 (SAXISCCTDATA_IN[144], SAXISCCTDATA[144]);
  buf B_SAXISCCTDATA145 (SAXISCCTDATA_IN[145], SAXISCCTDATA[145]);
  buf B_SAXISCCTDATA146 (SAXISCCTDATA_IN[146], SAXISCCTDATA[146]);
  buf B_SAXISCCTDATA147 (SAXISCCTDATA_IN[147], SAXISCCTDATA[147]);
  buf B_SAXISCCTDATA148 (SAXISCCTDATA_IN[148], SAXISCCTDATA[148]);
  buf B_SAXISCCTDATA149 (SAXISCCTDATA_IN[149], SAXISCCTDATA[149]);
  buf B_SAXISCCTDATA15 (SAXISCCTDATA_IN[15], SAXISCCTDATA[15]);
  buf B_SAXISCCTDATA150 (SAXISCCTDATA_IN[150], SAXISCCTDATA[150]);
  buf B_SAXISCCTDATA151 (SAXISCCTDATA_IN[151], SAXISCCTDATA[151]);
  buf B_SAXISCCTDATA152 (SAXISCCTDATA_IN[152], SAXISCCTDATA[152]);
  buf B_SAXISCCTDATA153 (SAXISCCTDATA_IN[153], SAXISCCTDATA[153]);
  buf B_SAXISCCTDATA154 (SAXISCCTDATA_IN[154], SAXISCCTDATA[154]);
  buf B_SAXISCCTDATA155 (SAXISCCTDATA_IN[155], SAXISCCTDATA[155]);
  buf B_SAXISCCTDATA156 (SAXISCCTDATA_IN[156], SAXISCCTDATA[156]);
  buf B_SAXISCCTDATA157 (SAXISCCTDATA_IN[157], SAXISCCTDATA[157]);
  buf B_SAXISCCTDATA158 (SAXISCCTDATA_IN[158], SAXISCCTDATA[158]);
  buf B_SAXISCCTDATA159 (SAXISCCTDATA_IN[159], SAXISCCTDATA[159]);
  buf B_SAXISCCTDATA16 (SAXISCCTDATA_IN[16], SAXISCCTDATA[16]);
  buf B_SAXISCCTDATA160 (SAXISCCTDATA_IN[160], SAXISCCTDATA[160]);
  buf B_SAXISCCTDATA161 (SAXISCCTDATA_IN[161], SAXISCCTDATA[161]);
  buf B_SAXISCCTDATA162 (SAXISCCTDATA_IN[162], SAXISCCTDATA[162]);
  buf B_SAXISCCTDATA163 (SAXISCCTDATA_IN[163], SAXISCCTDATA[163]);
  buf B_SAXISCCTDATA164 (SAXISCCTDATA_IN[164], SAXISCCTDATA[164]);
  buf B_SAXISCCTDATA165 (SAXISCCTDATA_IN[165], SAXISCCTDATA[165]);
  buf B_SAXISCCTDATA166 (SAXISCCTDATA_IN[166], SAXISCCTDATA[166]);
  buf B_SAXISCCTDATA167 (SAXISCCTDATA_IN[167], SAXISCCTDATA[167]);
  buf B_SAXISCCTDATA168 (SAXISCCTDATA_IN[168], SAXISCCTDATA[168]);
  buf B_SAXISCCTDATA169 (SAXISCCTDATA_IN[169], SAXISCCTDATA[169]);
  buf B_SAXISCCTDATA17 (SAXISCCTDATA_IN[17], SAXISCCTDATA[17]);
  buf B_SAXISCCTDATA170 (SAXISCCTDATA_IN[170], SAXISCCTDATA[170]);
  buf B_SAXISCCTDATA171 (SAXISCCTDATA_IN[171], SAXISCCTDATA[171]);
  buf B_SAXISCCTDATA172 (SAXISCCTDATA_IN[172], SAXISCCTDATA[172]);
  buf B_SAXISCCTDATA173 (SAXISCCTDATA_IN[173], SAXISCCTDATA[173]);
  buf B_SAXISCCTDATA174 (SAXISCCTDATA_IN[174], SAXISCCTDATA[174]);
  buf B_SAXISCCTDATA175 (SAXISCCTDATA_IN[175], SAXISCCTDATA[175]);
  buf B_SAXISCCTDATA176 (SAXISCCTDATA_IN[176], SAXISCCTDATA[176]);
  buf B_SAXISCCTDATA177 (SAXISCCTDATA_IN[177], SAXISCCTDATA[177]);
  buf B_SAXISCCTDATA178 (SAXISCCTDATA_IN[178], SAXISCCTDATA[178]);
  buf B_SAXISCCTDATA179 (SAXISCCTDATA_IN[179], SAXISCCTDATA[179]);
  buf B_SAXISCCTDATA18 (SAXISCCTDATA_IN[18], SAXISCCTDATA[18]);
  buf B_SAXISCCTDATA180 (SAXISCCTDATA_IN[180], SAXISCCTDATA[180]);
  buf B_SAXISCCTDATA181 (SAXISCCTDATA_IN[181], SAXISCCTDATA[181]);
  buf B_SAXISCCTDATA182 (SAXISCCTDATA_IN[182], SAXISCCTDATA[182]);
  buf B_SAXISCCTDATA183 (SAXISCCTDATA_IN[183], SAXISCCTDATA[183]);
  buf B_SAXISCCTDATA184 (SAXISCCTDATA_IN[184], SAXISCCTDATA[184]);
  buf B_SAXISCCTDATA185 (SAXISCCTDATA_IN[185], SAXISCCTDATA[185]);
  buf B_SAXISCCTDATA186 (SAXISCCTDATA_IN[186], SAXISCCTDATA[186]);
  buf B_SAXISCCTDATA187 (SAXISCCTDATA_IN[187], SAXISCCTDATA[187]);
  buf B_SAXISCCTDATA188 (SAXISCCTDATA_IN[188], SAXISCCTDATA[188]);
  buf B_SAXISCCTDATA189 (SAXISCCTDATA_IN[189], SAXISCCTDATA[189]);
  buf B_SAXISCCTDATA19 (SAXISCCTDATA_IN[19], SAXISCCTDATA[19]);
  buf B_SAXISCCTDATA190 (SAXISCCTDATA_IN[190], SAXISCCTDATA[190]);
  buf B_SAXISCCTDATA191 (SAXISCCTDATA_IN[191], SAXISCCTDATA[191]);
  buf B_SAXISCCTDATA192 (SAXISCCTDATA_IN[192], SAXISCCTDATA[192]);
  buf B_SAXISCCTDATA193 (SAXISCCTDATA_IN[193], SAXISCCTDATA[193]);
  buf B_SAXISCCTDATA194 (SAXISCCTDATA_IN[194], SAXISCCTDATA[194]);
  buf B_SAXISCCTDATA195 (SAXISCCTDATA_IN[195], SAXISCCTDATA[195]);
  buf B_SAXISCCTDATA196 (SAXISCCTDATA_IN[196], SAXISCCTDATA[196]);
  buf B_SAXISCCTDATA197 (SAXISCCTDATA_IN[197], SAXISCCTDATA[197]);
  buf B_SAXISCCTDATA198 (SAXISCCTDATA_IN[198], SAXISCCTDATA[198]);
  buf B_SAXISCCTDATA199 (SAXISCCTDATA_IN[199], SAXISCCTDATA[199]);
  buf B_SAXISCCTDATA2 (SAXISCCTDATA_IN[2], SAXISCCTDATA[2]);
  buf B_SAXISCCTDATA20 (SAXISCCTDATA_IN[20], SAXISCCTDATA[20]);
  buf B_SAXISCCTDATA200 (SAXISCCTDATA_IN[200], SAXISCCTDATA[200]);
  buf B_SAXISCCTDATA201 (SAXISCCTDATA_IN[201], SAXISCCTDATA[201]);
  buf B_SAXISCCTDATA202 (SAXISCCTDATA_IN[202], SAXISCCTDATA[202]);
  buf B_SAXISCCTDATA203 (SAXISCCTDATA_IN[203], SAXISCCTDATA[203]);
  buf B_SAXISCCTDATA204 (SAXISCCTDATA_IN[204], SAXISCCTDATA[204]);
  buf B_SAXISCCTDATA205 (SAXISCCTDATA_IN[205], SAXISCCTDATA[205]);
  buf B_SAXISCCTDATA206 (SAXISCCTDATA_IN[206], SAXISCCTDATA[206]);
  buf B_SAXISCCTDATA207 (SAXISCCTDATA_IN[207], SAXISCCTDATA[207]);
  buf B_SAXISCCTDATA208 (SAXISCCTDATA_IN[208], SAXISCCTDATA[208]);
  buf B_SAXISCCTDATA209 (SAXISCCTDATA_IN[209], SAXISCCTDATA[209]);
  buf B_SAXISCCTDATA21 (SAXISCCTDATA_IN[21], SAXISCCTDATA[21]);
  buf B_SAXISCCTDATA210 (SAXISCCTDATA_IN[210], SAXISCCTDATA[210]);
  buf B_SAXISCCTDATA211 (SAXISCCTDATA_IN[211], SAXISCCTDATA[211]);
  buf B_SAXISCCTDATA212 (SAXISCCTDATA_IN[212], SAXISCCTDATA[212]);
  buf B_SAXISCCTDATA213 (SAXISCCTDATA_IN[213], SAXISCCTDATA[213]);
  buf B_SAXISCCTDATA214 (SAXISCCTDATA_IN[214], SAXISCCTDATA[214]);
  buf B_SAXISCCTDATA215 (SAXISCCTDATA_IN[215], SAXISCCTDATA[215]);
  buf B_SAXISCCTDATA216 (SAXISCCTDATA_IN[216], SAXISCCTDATA[216]);
  buf B_SAXISCCTDATA217 (SAXISCCTDATA_IN[217], SAXISCCTDATA[217]);
  buf B_SAXISCCTDATA218 (SAXISCCTDATA_IN[218], SAXISCCTDATA[218]);
  buf B_SAXISCCTDATA219 (SAXISCCTDATA_IN[219], SAXISCCTDATA[219]);
  buf B_SAXISCCTDATA22 (SAXISCCTDATA_IN[22], SAXISCCTDATA[22]);
  buf B_SAXISCCTDATA220 (SAXISCCTDATA_IN[220], SAXISCCTDATA[220]);
  buf B_SAXISCCTDATA221 (SAXISCCTDATA_IN[221], SAXISCCTDATA[221]);
  buf B_SAXISCCTDATA222 (SAXISCCTDATA_IN[222], SAXISCCTDATA[222]);
  buf B_SAXISCCTDATA223 (SAXISCCTDATA_IN[223], SAXISCCTDATA[223]);
  buf B_SAXISCCTDATA224 (SAXISCCTDATA_IN[224], SAXISCCTDATA[224]);
  buf B_SAXISCCTDATA225 (SAXISCCTDATA_IN[225], SAXISCCTDATA[225]);
  buf B_SAXISCCTDATA226 (SAXISCCTDATA_IN[226], SAXISCCTDATA[226]);
  buf B_SAXISCCTDATA227 (SAXISCCTDATA_IN[227], SAXISCCTDATA[227]);
  buf B_SAXISCCTDATA228 (SAXISCCTDATA_IN[228], SAXISCCTDATA[228]);
  buf B_SAXISCCTDATA229 (SAXISCCTDATA_IN[229], SAXISCCTDATA[229]);
  buf B_SAXISCCTDATA23 (SAXISCCTDATA_IN[23], SAXISCCTDATA[23]);
  buf B_SAXISCCTDATA230 (SAXISCCTDATA_IN[230], SAXISCCTDATA[230]);
  buf B_SAXISCCTDATA231 (SAXISCCTDATA_IN[231], SAXISCCTDATA[231]);
  buf B_SAXISCCTDATA232 (SAXISCCTDATA_IN[232], SAXISCCTDATA[232]);
  buf B_SAXISCCTDATA233 (SAXISCCTDATA_IN[233], SAXISCCTDATA[233]);
  buf B_SAXISCCTDATA234 (SAXISCCTDATA_IN[234], SAXISCCTDATA[234]);
  buf B_SAXISCCTDATA235 (SAXISCCTDATA_IN[235], SAXISCCTDATA[235]);
  buf B_SAXISCCTDATA236 (SAXISCCTDATA_IN[236], SAXISCCTDATA[236]);
  buf B_SAXISCCTDATA237 (SAXISCCTDATA_IN[237], SAXISCCTDATA[237]);
  buf B_SAXISCCTDATA238 (SAXISCCTDATA_IN[238], SAXISCCTDATA[238]);
  buf B_SAXISCCTDATA239 (SAXISCCTDATA_IN[239], SAXISCCTDATA[239]);
  buf B_SAXISCCTDATA24 (SAXISCCTDATA_IN[24], SAXISCCTDATA[24]);
  buf B_SAXISCCTDATA240 (SAXISCCTDATA_IN[240], SAXISCCTDATA[240]);
  buf B_SAXISCCTDATA241 (SAXISCCTDATA_IN[241], SAXISCCTDATA[241]);
  buf B_SAXISCCTDATA242 (SAXISCCTDATA_IN[242], SAXISCCTDATA[242]);
  buf B_SAXISCCTDATA243 (SAXISCCTDATA_IN[243], SAXISCCTDATA[243]);
  buf B_SAXISCCTDATA244 (SAXISCCTDATA_IN[244], SAXISCCTDATA[244]);
  buf B_SAXISCCTDATA245 (SAXISCCTDATA_IN[245], SAXISCCTDATA[245]);
  buf B_SAXISCCTDATA246 (SAXISCCTDATA_IN[246], SAXISCCTDATA[246]);
  buf B_SAXISCCTDATA247 (SAXISCCTDATA_IN[247], SAXISCCTDATA[247]);
  buf B_SAXISCCTDATA248 (SAXISCCTDATA_IN[248], SAXISCCTDATA[248]);
  buf B_SAXISCCTDATA249 (SAXISCCTDATA_IN[249], SAXISCCTDATA[249]);
  buf B_SAXISCCTDATA25 (SAXISCCTDATA_IN[25], SAXISCCTDATA[25]);
  buf B_SAXISCCTDATA250 (SAXISCCTDATA_IN[250], SAXISCCTDATA[250]);
  buf B_SAXISCCTDATA251 (SAXISCCTDATA_IN[251], SAXISCCTDATA[251]);
  buf B_SAXISCCTDATA252 (SAXISCCTDATA_IN[252], SAXISCCTDATA[252]);
  buf B_SAXISCCTDATA253 (SAXISCCTDATA_IN[253], SAXISCCTDATA[253]);
  buf B_SAXISCCTDATA254 (SAXISCCTDATA_IN[254], SAXISCCTDATA[254]);
  buf B_SAXISCCTDATA255 (SAXISCCTDATA_IN[255], SAXISCCTDATA[255]);
  buf B_SAXISCCTDATA26 (SAXISCCTDATA_IN[26], SAXISCCTDATA[26]);
  buf B_SAXISCCTDATA27 (SAXISCCTDATA_IN[27], SAXISCCTDATA[27]);
  buf B_SAXISCCTDATA28 (SAXISCCTDATA_IN[28], SAXISCCTDATA[28]);
  buf B_SAXISCCTDATA29 (SAXISCCTDATA_IN[29], SAXISCCTDATA[29]);
  buf B_SAXISCCTDATA3 (SAXISCCTDATA_IN[3], SAXISCCTDATA[3]);
  buf B_SAXISCCTDATA30 (SAXISCCTDATA_IN[30], SAXISCCTDATA[30]);
  buf B_SAXISCCTDATA31 (SAXISCCTDATA_IN[31], SAXISCCTDATA[31]);
  buf B_SAXISCCTDATA32 (SAXISCCTDATA_IN[32], SAXISCCTDATA[32]);
  buf B_SAXISCCTDATA33 (SAXISCCTDATA_IN[33], SAXISCCTDATA[33]);
  buf B_SAXISCCTDATA34 (SAXISCCTDATA_IN[34], SAXISCCTDATA[34]);
  buf B_SAXISCCTDATA35 (SAXISCCTDATA_IN[35], SAXISCCTDATA[35]);
  buf B_SAXISCCTDATA36 (SAXISCCTDATA_IN[36], SAXISCCTDATA[36]);
  buf B_SAXISCCTDATA37 (SAXISCCTDATA_IN[37], SAXISCCTDATA[37]);
  buf B_SAXISCCTDATA38 (SAXISCCTDATA_IN[38], SAXISCCTDATA[38]);
  buf B_SAXISCCTDATA39 (SAXISCCTDATA_IN[39], SAXISCCTDATA[39]);
  buf B_SAXISCCTDATA4 (SAXISCCTDATA_IN[4], SAXISCCTDATA[4]);
  buf B_SAXISCCTDATA40 (SAXISCCTDATA_IN[40], SAXISCCTDATA[40]);
  buf B_SAXISCCTDATA41 (SAXISCCTDATA_IN[41], SAXISCCTDATA[41]);
  buf B_SAXISCCTDATA42 (SAXISCCTDATA_IN[42], SAXISCCTDATA[42]);
  buf B_SAXISCCTDATA43 (SAXISCCTDATA_IN[43], SAXISCCTDATA[43]);
  buf B_SAXISCCTDATA44 (SAXISCCTDATA_IN[44], SAXISCCTDATA[44]);
  buf B_SAXISCCTDATA45 (SAXISCCTDATA_IN[45], SAXISCCTDATA[45]);
  buf B_SAXISCCTDATA46 (SAXISCCTDATA_IN[46], SAXISCCTDATA[46]);
  buf B_SAXISCCTDATA47 (SAXISCCTDATA_IN[47], SAXISCCTDATA[47]);
  buf B_SAXISCCTDATA48 (SAXISCCTDATA_IN[48], SAXISCCTDATA[48]);
  buf B_SAXISCCTDATA49 (SAXISCCTDATA_IN[49], SAXISCCTDATA[49]);
  buf B_SAXISCCTDATA5 (SAXISCCTDATA_IN[5], SAXISCCTDATA[5]);
  buf B_SAXISCCTDATA50 (SAXISCCTDATA_IN[50], SAXISCCTDATA[50]);
  buf B_SAXISCCTDATA51 (SAXISCCTDATA_IN[51], SAXISCCTDATA[51]);
  buf B_SAXISCCTDATA52 (SAXISCCTDATA_IN[52], SAXISCCTDATA[52]);
  buf B_SAXISCCTDATA53 (SAXISCCTDATA_IN[53], SAXISCCTDATA[53]);
  buf B_SAXISCCTDATA54 (SAXISCCTDATA_IN[54], SAXISCCTDATA[54]);
  buf B_SAXISCCTDATA55 (SAXISCCTDATA_IN[55], SAXISCCTDATA[55]);
  buf B_SAXISCCTDATA56 (SAXISCCTDATA_IN[56], SAXISCCTDATA[56]);
  buf B_SAXISCCTDATA57 (SAXISCCTDATA_IN[57], SAXISCCTDATA[57]);
  buf B_SAXISCCTDATA58 (SAXISCCTDATA_IN[58], SAXISCCTDATA[58]);
  buf B_SAXISCCTDATA59 (SAXISCCTDATA_IN[59], SAXISCCTDATA[59]);
  buf B_SAXISCCTDATA6 (SAXISCCTDATA_IN[6], SAXISCCTDATA[6]);
  buf B_SAXISCCTDATA60 (SAXISCCTDATA_IN[60], SAXISCCTDATA[60]);
  buf B_SAXISCCTDATA61 (SAXISCCTDATA_IN[61], SAXISCCTDATA[61]);
  buf B_SAXISCCTDATA62 (SAXISCCTDATA_IN[62], SAXISCCTDATA[62]);
  buf B_SAXISCCTDATA63 (SAXISCCTDATA_IN[63], SAXISCCTDATA[63]);
  buf B_SAXISCCTDATA64 (SAXISCCTDATA_IN[64], SAXISCCTDATA[64]);
  buf B_SAXISCCTDATA65 (SAXISCCTDATA_IN[65], SAXISCCTDATA[65]);
  buf B_SAXISCCTDATA66 (SAXISCCTDATA_IN[66], SAXISCCTDATA[66]);
  buf B_SAXISCCTDATA67 (SAXISCCTDATA_IN[67], SAXISCCTDATA[67]);
  buf B_SAXISCCTDATA68 (SAXISCCTDATA_IN[68], SAXISCCTDATA[68]);
  buf B_SAXISCCTDATA69 (SAXISCCTDATA_IN[69], SAXISCCTDATA[69]);
  buf B_SAXISCCTDATA7 (SAXISCCTDATA_IN[7], SAXISCCTDATA[7]);
  buf B_SAXISCCTDATA70 (SAXISCCTDATA_IN[70], SAXISCCTDATA[70]);
  buf B_SAXISCCTDATA71 (SAXISCCTDATA_IN[71], SAXISCCTDATA[71]);
  buf B_SAXISCCTDATA72 (SAXISCCTDATA_IN[72], SAXISCCTDATA[72]);
  buf B_SAXISCCTDATA73 (SAXISCCTDATA_IN[73], SAXISCCTDATA[73]);
  buf B_SAXISCCTDATA74 (SAXISCCTDATA_IN[74], SAXISCCTDATA[74]);
  buf B_SAXISCCTDATA75 (SAXISCCTDATA_IN[75], SAXISCCTDATA[75]);
  buf B_SAXISCCTDATA76 (SAXISCCTDATA_IN[76], SAXISCCTDATA[76]);
  buf B_SAXISCCTDATA77 (SAXISCCTDATA_IN[77], SAXISCCTDATA[77]);
  buf B_SAXISCCTDATA78 (SAXISCCTDATA_IN[78], SAXISCCTDATA[78]);
  buf B_SAXISCCTDATA79 (SAXISCCTDATA_IN[79], SAXISCCTDATA[79]);
  buf B_SAXISCCTDATA8 (SAXISCCTDATA_IN[8], SAXISCCTDATA[8]);
  buf B_SAXISCCTDATA80 (SAXISCCTDATA_IN[80], SAXISCCTDATA[80]);
  buf B_SAXISCCTDATA81 (SAXISCCTDATA_IN[81], SAXISCCTDATA[81]);
  buf B_SAXISCCTDATA82 (SAXISCCTDATA_IN[82], SAXISCCTDATA[82]);
  buf B_SAXISCCTDATA83 (SAXISCCTDATA_IN[83], SAXISCCTDATA[83]);
  buf B_SAXISCCTDATA84 (SAXISCCTDATA_IN[84], SAXISCCTDATA[84]);
  buf B_SAXISCCTDATA85 (SAXISCCTDATA_IN[85], SAXISCCTDATA[85]);
  buf B_SAXISCCTDATA86 (SAXISCCTDATA_IN[86], SAXISCCTDATA[86]);
  buf B_SAXISCCTDATA87 (SAXISCCTDATA_IN[87], SAXISCCTDATA[87]);
  buf B_SAXISCCTDATA88 (SAXISCCTDATA_IN[88], SAXISCCTDATA[88]);
  buf B_SAXISCCTDATA89 (SAXISCCTDATA_IN[89], SAXISCCTDATA[89]);
  buf B_SAXISCCTDATA9 (SAXISCCTDATA_IN[9], SAXISCCTDATA[9]);
  buf B_SAXISCCTDATA90 (SAXISCCTDATA_IN[90], SAXISCCTDATA[90]);
  buf B_SAXISCCTDATA91 (SAXISCCTDATA_IN[91], SAXISCCTDATA[91]);
  buf B_SAXISCCTDATA92 (SAXISCCTDATA_IN[92], SAXISCCTDATA[92]);
  buf B_SAXISCCTDATA93 (SAXISCCTDATA_IN[93], SAXISCCTDATA[93]);
  buf B_SAXISCCTDATA94 (SAXISCCTDATA_IN[94], SAXISCCTDATA[94]);
  buf B_SAXISCCTDATA95 (SAXISCCTDATA_IN[95], SAXISCCTDATA[95]);
  buf B_SAXISCCTDATA96 (SAXISCCTDATA_IN[96], SAXISCCTDATA[96]);
  buf B_SAXISCCTDATA97 (SAXISCCTDATA_IN[97], SAXISCCTDATA[97]);
  buf B_SAXISCCTDATA98 (SAXISCCTDATA_IN[98], SAXISCCTDATA[98]);
  buf B_SAXISCCTDATA99 (SAXISCCTDATA_IN[99], SAXISCCTDATA[99]);
  buf B_SAXISCCTKEEP0 (SAXISCCTKEEP_IN[0], SAXISCCTKEEP[0]);
  buf B_SAXISCCTKEEP1 (SAXISCCTKEEP_IN[1], SAXISCCTKEEP[1]);
  buf B_SAXISCCTKEEP2 (SAXISCCTKEEP_IN[2], SAXISCCTKEEP[2]);
  buf B_SAXISCCTKEEP3 (SAXISCCTKEEP_IN[3], SAXISCCTKEEP[3]);
  buf B_SAXISCCTKEEP4 (SAXISCCTKEEP_IN[4], SAXISCCTKEEP[4]);
  buf B_SAXISCCTKEEP5 (SAXISCCTKEEP_IN[5], SAXISCCTKEEP[5]);
  buf B_SAXISCCTKEEP6 (SAXISCCTKEEP_IN[6], SAXISCCTKEEP[6]);
  buf B_SAXISCCTKEEP7 (SAXISCCTKEEP_IN[7], SAXISCCTKEEP[7]);
  buf B_SAXISCCTLAST (SAXISCCTLAST_IN, SAXISCCTLAST);
  buf B_SAXISCCTUSER0 (SAXISCCTUSER_IN[0], SAXISCCTUSER[0]);
  buf B_SAXISCCTUSER1 (SAXISCCTUSER_IN[1], SAXISCCTUSER[1]);
  buf B_SAXISCCTUSER10 (SAXISCCTUSER_IN[10], SAXISCCTUSER[10]);
  buf B_SAXISCCTUSER11 (SAXISCCTUSER_IN[11], SAXISCCTUSER[11]);
  buf B_SAXISCCTUSER12 (SAXISCCTUSER_IN[12], SAXISCCTUSER[12]);
  buf B_SAXISCCTUSER13 (SAXISCCTUSER_IN[13], SAXISCCTUSER[13]);
  buf B_SAXISCCTUSER14 (SAXISCCTUSER_IN[14], SAXISCCTUSER[14]);
  buf B_SAXISCCTUSER15 (SAXISCCTUSER_IN[15], SAXISCCTUSER[15]);
  buf B_SAXISCCTUSER16 (SAXISCCTUSER_IN[16], SAXISCCTUSER[16]);
  buf B_SAXISCCTUSER17 (SAXISCCTUSER_IN[17], SAXISCCTUSER[17]);
  buf B_SAXISCCTUSER18 (SAXISCCTUSER_IN[18], SAXISCCTUSER[18]);
  buf B_SAXISCCTUSER19 (SAXISCCTUSER_IN[19], SAXISCCTUSER[19]);
  buf B_SAXISCCTUSER2 (SAXISCCTUSER_IN[2], SAXISCCTUSER[2]);
  buf B_SAXISCCTUSER20 (SAXISCCTUSER_IN[20], SAXISCCTUSER[20]);
  buf B_SAXISCCTUSER21 (SAXISCCTUSER_IN[21], SAXISCCTUSER[21]);
  buf B_SAXISCCTUSER22 (SAXISCCTUSER_IN[22], SAXISCCTUSER[22]);
  buf B_SAXISCCTUSER23 (SAXISCCTUSER_IN[23], SAXISCCTUSER[23]);
  buf B_SAXISCCTUSER24 (SAXISCCTUSER_IN[24], SAXISCCTUSER[24]);
  buf B_SAXISCCTUSER25 (SAXISCCTUSER_IN[25], SAXISCCTUSER[25]);
  buf B_SAXISCCTUSER26 (SAXISCCTUSER_IN[26], SAXISCCTUSER[26]);
  buf B_SAXISCCTUSER27 (SAXISCCTUSER_IN[27], SAXISCCTUSER[27]);
  buf B_SAXISCCTUSER28 (SAXISCCTUSER_IN[28], SAXISCCTUSER[28]);
  buf B_SAXISCCTUSER29 (SAXISCCTUSER_IN[29], SAXISCCTUSER[29]);
  buf B_SAXISCCTUSER3 (SAXISCCTUSER_IN[3], SAXISCCTUSER[3]);
  buf B_SAXISCCTUSER30 (SAXISCCTUSER_IN[30], SAXISCCTUSER[30]);
  buf B_SAXISCCTUSER31 (SAXISCCTUSER_IN[31], SAXISCCTUSER[31]);
  buf B_SAXISCCTUSER32 (SAXISCCTUSER_IN[32], SAXISCCTUSER[32]);
  buf B_SAXISCCTUSER4 (SAXISCCTUSER_IN[4], SAXISCCTUSER[4]);
  buf B_SAXISCCTUSER5 (SAXISCCTUSER_IN[5], SAXISCCTUSER[5]);
  buf B_SAXISCCTUSER6 (SAXISCCTUSER_IN[6], SAXISCCTUSER[6]);
  buf B_SAXISCCTUSER7 (SAXISCCTUSER_IN[7], SAXISCCTUSER[7]);
  buf B_SAXISCCTUSER8 (SAXISCCTUSER_IN[8], SAXISCCTUSER[8]);
  buf B_SAXISCCTUSER9 (SAXISCCTUSER_IN[9], SAXISCCTUSER[9]);
  buf B_SAXISCCTVALID (SAXISCCTVALID_IN, SAXISCCTVALID);
  buf B_SAXISRQTDATA0 (SAXISRQTDATA_IN[0], SAXISRQTDATA[0]);
  buf B_SAXISRQTDATA1 (SAXISRQTDATA_IN[1], SAXISRQTDATA[1]);
  buf B_SAXISRQTDATA10 (SAXISRQTDATA_IN[10], SAXISRQTDATA[10]);
  buf B_SAXISRQTDATA100 (SAXISRQTDATA_IN[100], SAXISRQTDATA[100]);
  buf B_SAXISRQTDATA101 (SAXISRQTDATA_IN[101], SAXISRQTDATA[101]);
  buf B_SAXISRQTDATA102 (SAXISRQTDATA_IN[102], SAXISRQTDATA[102]);
  buf B_SAXISRQTDATA103 (SAXISRQTDATA_IN[103], SAXISRQTDATA[103]);
  buf B_SAXISRQTDATA104 (SAXISRQTDATA_IN[104], SAXISRQTDATA[104]);
  buf B_SAXISRQTDATA105 (SAXISRQTDATA_IN[105], SAXISRQTDATA[105]);
  buf B_SAXISRQTDATA106 (SAXISRQTDATA_IN[106], SAXISRQTDATA[106]);
  buf B_SAXISRQTDATA107 (SAXISRQTDATA_IN[107], SAXISRQTDATA[107]);
  buf B_SAXISRQTDATA108 (SAXISRQTDATA_IN[108], SAXISRQTDATA[108]);
  buf B_SAXISRQTDATA109 (SAXISRQTDATA_IN[109], SAXISRQTDATA[109]);
  buf B_SAXISRQTDATA11 (SAXISRQTDATA_IN[11], SAXISRQTDATA[11]);
  buf B_SAXISRQTDATA110 (SAXISRQTDATA_IN[110], SAXISRQTDATA[110]);
  buf B_SAXISRQTDATA111 (SAXISRQTDATA_IN[111], SAXISRQTDATA[111]);
  buf B_SAXISRQTDATA112 (SAXISRQTDATA_IN[112], SAXISRQTDATA[112]);
  buf B_SAXISRQTDATA113 (SAXISRQTDATA_IN[113], SAXISRQTDATA[113]);
  buf B_SAXISRQTDATA114 (SAXISRQTDATA_IN[114], SAXISRQTDATA[114]);
  buf B_SAXISRQTDATA115 (SAXISRQTDATA_IN[115], SAXISRQTDATA[115]);
  buf B_SAXISRQTDATA116 (SAXISRQTDATA_IN[116], SAXISRQTDATA[116]);
  buf B_SAXISRQTDATA117 (SAXISRQTDATA_IN[117], SAXISRQTDATA[117]);
  buf B_SAXISRQTDATA118 (SAXISRQTDATA_IN[118], SAXISRQTDATA[118]);
  buf B_SAXISRQTDATA119 (SAXISRQTDATA_IN[119], SAXISRQTDATA[119]);
  buf B_SAXISRQTDATA12 (SAXISRQTDATA_IN[12], SAXISRQTDATA[12]);
  buf B_SAXISRQTDATA120 (SAXISRQTDATA_IN[120], SAXISRQTDATA[120]);
  buf B_SAXISRQTDATA121 (SAXISRQTDATA_IN[121], SAXISRQTDATA[121]);
  buf B_SAXISRQTDATA122 (SAXISRQTDATA_IN[122], SAXISRQTDATA[122]);
  buf B_SAXISRQTDATA123 (SAXISRQTDATA_IN[123], SAXISRQTDATA[123]);
  buf B_SAXISRQTDATA124 (SAXISRQTDATA_IN[124], SAXISRQTDATA[124]);
  buf B_SAXISRQTDATA125 (SAXISRQTDATA_IN[125], SAXISRQTDATA[125]);
  buf B_SAXISRQTDATA126 (SAXISRQTDATA_IN[126], SAXISRQTDATA[126]);
  buf B_SAXISRQTDATA127 (SAXISRQTDATA_IN[127], SAXISRQTDATA[127]);
  buf B_SAXISRQTDATA128 (SAXISRQTDATA_IN[128], SAXISRQTDATA[128]);
  buf B_SAXISRQTDATA129 (SAXISRQTDATA_IN[129], SAXISRQTDATA[129]);
  buf B_SAXISRQTDATA13 (SAXISRQTDATA_IN[13], SAXISRQTDATA[13]);
  buf B_SAXISRQTDATA130 (SAXISRQTDATA_IN[130], SAXISRQTDATA[130]);
  buf B_SAXISRQTDATA131 (SAXISRQTDATA_IN[131], SAXISRQTDATA[131]);
  buf B_SAXISRQTDATA132 (SAXISRQTDATA_IN[132], SAXISRQTDATA[132]);
  buf B_SAXISRQTDATA133 (SAXISRQTDATA_IN[133], SAXISRQTDATA[133]);
  buf B_SAXISRQTDATA134 (SAXISRQTDATA_IN[134], SAXISRQTDATA[134]);
  buf B_SAXISRQTDATA135 (SAXISRQTDATA_IN[135], SAXISRQTDATA[135]);
  buf B_SAXISRQTDATA136 (SAXISRQTDATA_IN[136], SAXISRQTDATA[136]);
  buf B_SAXISRQTDATA137 (SAXISRQTDATA_IN[137], SAXISRQTDATA[137]);
  buf B_SAXISRQTDATA138 (SAXISRQTDATA_IN[138], SAXISRQTDATA[138]);
  buf B_SAXISRQTDATA139 (SAXISRQTDATA_IN[139], SAXISRQTDATA[139]);
  buf B_SAXISRQTDATA14 (SAXISRQTDATA_IN[14], SAXISRQTDATA[14]);
  buf B_SAXISRQTDATA140 (SAXISRQTDATA_IN[140], SAXISRQTDATA[140]);
  buf B_SAXISRQTDATA141 (SAXISRQTDATA_IN[141], SAXISRQTDATA[141]);
  buf B_SAXISRQTDATA142 (SAXISRQTDATA_IN[142], SAXISRQTDATA[142]);
  buf B_SAXISRQTDATA143 (SAXISRQTDATA_IN[143], SAXISRQTDATA[143]);
  buf B_SAXISRQTDATA144 (SAXISRQTDATA_IN[144], SAXISRQTDATA[144]);
  buf B_SAXISRQTDATA145 (SAXISRQTDATA_IN[145], SAXISRQTDATA[145]);
  buf B_SAXISRQTDATA146 (SAXISRQTDATA_IN[146], SAXISRQTDATA[146]);
  buf B_SAXISRQTDATA147 (SAXISRQTDATA_IN[147], SAXISRQTDATA[147]);
  buf B_SAXISRQTDATA148 (SAXISRQTDATA_IN[148], SAXISRQTDATA[148]);
  buf B_SAXISRQTDATA149 (SAXISRQTDATA_IN[149], SAXISRQTDATA[149]);
  buf B_SAXISRQTDATA15 (SAXISRQTDATA_IN[15], SAXISRQTDATA[15]);
  buf B_SAXISRQTDATA150 (SAXISRQTDATA_IN[150], SAXISRQTDATA[150]);
  buf B_SAXISRQTDATA151 (SAXISRQTDATA_IN[151], SAXISRQTDATA[151]);
  buf B_SAXISRQTDATA152 (SAXISRQTDATA_IN[152], SAXISRQTDATA[152]);
  buf B_SAXISRQTDATA153 (SAXISRQTDATA_IN[153], SAXISRQTDATA[153]);
  buf B_SAXISRQTDATA154 (SAXISRQTDATA_IN[154], SAXISRQTDATA[154]);
  buf B_SAXISRQTDATA155 (SAXISRQTDATA_IN[155], SAXISRQTDATA[155]);
  buf B_SAXISRQTDATA156 (SAXISRQTDATA_IN[156], SAXISRQTDATA[156]);
  buf B_SAXISRQTDATA157 (SAXISRQTDATA_IN[157], SAXISRQTDATA[157]);
  buf B_SAXISRQTDATA158 (SAXISRQTDATA_IN[158], SAXISRQTDATA[158]);
  buf B_SAXISRQTDATA159 (SAXISRQTDATA_IN[159], SAXISRQTDATA[159]);
  buf B_SAXISRQTDATA16 (SAXISRQTDATA_IN[16], SAXISRQTDATA[16]);
  buf B_SAXISRQTDATA160 (SAXISRQTDATA_IN[160], SAXISRQTDATA[160]);
  buf B_SAXISRQTDATA161 (SAXISRQTDATA_IN[161], SAXISRQTDATA[161]);
  buf B_SAXISRQTDATA162 (SAXISRQTDATA_IN[162], SAXISRQTDATA[162]);
  buf B_SAXISRQTDATA163 (SAXISRQTDATA_IN[163], SAXISRQTDATA[163]);
  buf B_SAXISRQTDATA164 (SAXISRQTDATA_IN[164], SAXISRQTDATA[164]);
  buf B_SAXISRQTDATA165 (SAXISRQTDATA_IN[165], SAXISRQTDATA[165]);
  buf B_SAXISRQTDATA166 (SAXISRQTDATA_IN[166], SAXISRQTDATA[166]);
  buf B_SAXISRQTDATA167 (SAXISRQTDATA_IN[167], SAXISRQTDATA[167]);
  buf B_SAXISRQTDATA168 (SAXISRQTDATA_IN[168], SAXISRQTDATA[168]);
  buf B_SAXISRQTDATA169 (SAXISRQTDATA_IN[169], SAXISRQTDATA[169]);
  buf B_SAXISRQTDATA17 (SAXISRQTDATA_IN[17], SAXISRQTDATA[17]);
  buf B_SAXISRQTDATA170 (SAXISRQTDATA_IN[170], SAXISRQTDATA[170]);
  buf B_SAXISRQTDATA171 (SAXISRQTDATA_IN[171], SAXISRQTDATA[171]);
  buf B_SAXISRQTDATA172 (SAXISRQTDATA_IN[172], SAXISRQTDATA[172]);
  buf B_SAXISRQTDATA173 (SAXISRQTDATA_IN[173], SAXISRQTDATA[173]);
  buf B_SAXISRQTDATA174 (SAXISRQTDATA_IN[174], SAXISRQTDATA[174]);
  buf B_SAXISRQTDATA175 (SAXISRQTDATA_IN[175], SAXISRQTDATA[175]);
  buf B_SAXISRQTDATA176 (SAXISRQTDATA_IN[176], SAXISRQTDATA[176]);
  buf B_SAXISRQTDATA177 (SAXISRQTDATA_IN[177], SAXISRQTDATA[177]);
  buf B_SAXISRQTDATA178 (SAXISRQTDATA_IN[178], SAXISRQTDATA[178]);
  buf B_SAXISRQTDATA179 (SAXISRQTDATA_IN[179], SAXISRQTDATA[179]);
  buf B_SAXISRQTDATA18 (SAXISRQTDATA_IN[18], SAXISRQTDATA[18]);
  buf B_SAXISRQTDATA180 (SAXISRQTDATA_IN[180], SAXISRQTDATA[180]);
  buf B_SAXISRQTDATA181 (SAXISRQTDATA_IN[181], SAXISRQTDATA[181]);
  buf B_SAXISRQTDATA182 (SAXISRQTDATA_IN[182], SAXISRQTDATA[182]);
  buf B_SAXISRQTDATA183 (SAXISRQTDATA_IN[183], SAXISRQTDATA[183]);
  buf B_SAXISRQTDATA184 (SAXISRQTDATA_IN[184], SAXISRQTDATA[184]);
  buf B_SAXISRQTDATA185 (SAXISRQTDATA_IN[185], SAXISRQTDATA[185]);
  buf B_SAXISRQTDATA186 (SAXISRQTDATA_IN[186], SAXISRQTDATA[186]);
  buf B_SAXISRQTDATA187 (SAXISRQTDATA_IN[187], SAXISRQTDATA[187]);
  buf B_SAXISRQTDATA188 (SAXISRQTDATA_IN[188], SAXISRQTDATA[188]);
  buf B_SAXISRQTDATA189 (SAXISRQTDATA_IN[189], SAXISRQTDATA[189]);
  buf B_SAXISRQTDATA19 (SAXISRQTDATA_IN[19], SAXISRQTDATA[19]);
  buf B_SAXISRQTDATA190 (SAXISRQTDATA_IN[190], SAXISRQTDATA[190]);
  buf B_SAXISRQTDATA191 (SAXISRQTDATA_IN[191], SAXISRQTDATA[191]);
  buf B_SAXISRQTDATA192 (SAXISRQTDATA_IN[192], SAXISRQTDATA[192]);
  buf B_SAXISRQTDATA193 (SAXISRQTDATA_IN[193], SAXISRQTDATA[193]);
  buf B_SAXISRQTDATA194 (SAXISRQTDATA_IN[194], SAXISRQTDATA[194]);
  buf B_SAXISRQTDATA195 (SAXISRQTDATA_IN[195], SAXISRQTDATA[195]);
  buf B_SAXISRQTDATA196 (SAXISRQTDATA_IN[196], SAXISRQTDATA[196]);
  buf B_SAXISRQTDATA197 (SAXISRQTDATA_IN[197], SAXISRQTDATA[197]);
  buf B_SAXISRQTDATA198 (SAXISRQTDATA_IN[198], SAXISRQTDATA[198]);
  buf B_SAXISRQTDATA199 (SAXISRQTDATA_IN[199], SAXISRQTDATA[199]);
  buf B_SAXISRQTDATA2 (SAXISRQTDATA_IN[2], SAXISRQTDATA[2]);
  buf B_SAXISRQTDATA20 (SAXISRQTDATA_IN[20], SAXISRQTDATA[20]);
  buf B_SAXISRQTDATA200 (SAXISRQTDATA_IN[200], SAXISRQTDATA[200]);
  buf B_SAXISRQTDATA201 (SAXISRQTDATA_IN[201], SAXISRQTDATA[201]);
  buf B_SAXISRQTDATA202 (SAXISRQTDATA_IN[202], SAXISRQTDATA[202]);
  buf B_SAXISRQTDATA203 (SAXISRQTDATA_IN[203], SAXISRQTDATA[203]);
  buf B_SAXISRQTDATA204 (SAXISRQTDATA_IN[204], SAXISRQTDATA[204]);
  buf B_SAXISRQTDATA205 (SAXISRQTDATA_IN[205], SAXISRQTDATA[205]);
  buf B_SAXISRQTDATA206 (SAXISRQTDATA_IN[206], SAXISRQTDATA[206]);
  buf B_SAXISRQTDATA207 (SAXISRQTDATA_IN[207], SAXISRQTDATA[207]);
  buf B_SAXISRQTDATA208 (SAXISRQTDATA_IN[208], SAXISRQTDATA[208]);
  buf B_SAXISRQTDATA209 (SAXISRQTDATA_IN[209], SAXISRQTDATA[209]);
  buf B_SAXISRQTDATA21 (SAXISRQTDATA_IN[21], SAXISRQTDATA[21]);
  buf B_SAXISRQTDATA210 (SAXISRQTDATA_IN[210], SAXISRQTDATA[210]);
  buf B_SAXISRQTDATA211 (SAXISRQTDATA_IN[211], SAXISRQTDATA[211]);
  buf B_SAXISRQTDATA212 (SAXISRQTDATA_IN[212], SAXISRQTDATA[212]);
  buf B_SAXISRQTDATA213 (SAXISRQTDATA_IN[213], SAXISRQTDATA[213]);
  buf B_SAXISRQTDATA214 (SAXISRQTDATA_IN[214], SAXISRQTDATA[214]);
  buf B_SAXISRQTDATA215 (SAXISRQTDATA_IN[215], SAXISRQTDATA[215]);
  buf B_SAXISRQTDATA216 (SAXISRQTDATA_IN[216], SAXISRQTDATA[216]);
  buf B_SAXISRQTDATA217 (SAXISRQTDATA_IN[217], SAXISRQTDATA[217]);
  buf B_SAXISRQTDATA218 (SAXISRQTDATA_IN[218], SAXISRQTDATA[218]);
  buf B_SAXISRQTDATA219 (SAXISRQTDATA_IN[219], SAXISRQTDATA[219]);
  buf B_SAXISRQTDATA22 (SAXISRQTDATA_IN[22], SAXISRQTDATA[22]);
  buf B_SAXISRQTDATA220 (SAXISRQTDATA_IN[220], SAXISRQTDATA[220]);
  buf B_SAXISRQTDATA221 (SAXISRQTDATA_IN[221], SAXISRQTDATA[221]);
  buf B_SAXISRQTDATA222 (SAXISRQTDATA_IN[222], SAXISRQTDATA[222]);
  buf B_SAXISRQTDATA223 (SAXISRQTDATA_IN[223], SAXISRQTDATA[223]);
  buf B_SAXISRQTDATA224 (SAXISRQTDATA_IN[224], SAXISRQTDATA[224]);
  buf B_SAXISRQTDATA225 (SAXISRQTDATA_IN[225], SAXISRQTDATA[225]);
  buf B_SAXISRQTDATA226 (SAXISRQTDATA_IN[226], SAXISRQTDATA[226]);
  buf B_SAXISRQTDATA227 (SAXISRQTDATA_IN[227], SAXISRQTDATA[227]);
  buf B_SAXISRQTDATA228 (SAXISRQTDATA_IN[228], SAXISRQTDATA[228]);
  buf B_SAXISRQTDATA229 (SAXISRQTDATA_IN[229], SAXISRQTDATA[229]);
  buf B_SAXISRQTDATA23 (SAXISRQTDATA_IN[23], SAXISRQTDATA[23]);
  buf B_SAXISRQTDATA230 (SAXISRQTDATA_IN[230], SAXISRQTDATA[230]);
  buf B_SAXISRQTDATA231 (SAXISRQTDATA_IN[231], SAXISRQTDATA[231]);
  buf B_SAXISRQTDATA232 (SAXISRQTDATA_IN[232], SAXISRQTDATA[232]);
  buf B_SAXISRQTDATA233 (SAXISRQTDATA_IN[233], SAXISRQTDATA[233]);
  buf B_SAXISRQTDATA234 (SAXISRQTDATA_IN[234], SAXISRQTDATA[234]);
  buf B_SAXISRQTDATA235 (SAXISRQTDATA_IN[235], SAXISRQTDATA[235]);
  buf B_SAXISRQTDATA236 (SAXISRQTDATA_IN[236], SAXISRQTDATA[236]);
  buf B_SAXISRQTDATA237 (SAXISRQTDATA_IN[237], SAXISRQTDATA[237]);
  buf B_SAXISRQTDATA238 (SAXISRQTDATA_IN[238], SAXISRQTDATA[238]);
  buf B_SAXISRQTDATA239 (SAXISRQTDATA_IN[239], SAXISRQTDATA[239]);
  buf B_SAXISRQTDATA24 (SAXISRQTDATA_IN[24], SAXISRQTDATA[24]);
  buf B_SAXISRQTDATA240 (SAXISRQTDATA_IN[240], SAXISRQTDATA[240]);
  buf B_SAXISRQTDATA241 (SAXISRQTDATA_IN[241], SAXISRQTDATA[241]);
  buf B_SAXISRQTDATA242 (SAXISRQTDATA_IN[242], SAXISRQTDATA[242]);
  buf B_SAXISRQTDATA243 (SAXISRQTDATA_IN[243], SAXISRQTDATA[243]);
  buf B_SAXISRQTDATA244 (SAXISRQTDATA_IN[244], SAXISRQTDATA[244]);
  buf B_SAXISRQTDATA245 (SAXISRQTDATA_IN[245], SAXISRQTDATA[245]);
  buf B_SAXISRQTDATA246 (SAXISRQTDATA_IN[246], SAXISRQTDATA[246]);
  buf B_SAXISRQTDATA247 (SAXISRQTDATA_IN[247], SAXISRQTDATA[247]);
  buf B_SAXISRQTDATA248 (SAXISRQTDATA_IN[248], SAXISRQTDATA[248]);
  buf B_SAXISRQTDATA249 (SAXISRQTDATA_IN[249], SAXISRQTDATA[249]);
  buf B_SAXISRQTDATA25 (SAXISRQTDATA_IN[25], SAXISRQTDATA[25]);
  buf B_SAXISRQTDATA250 (SAXISRQTDATA_IN[250], SAXISRQTDATA[250]);
  buf B_SAXISRQTDATA251 (SAXISRQTDATA_IN[251], SAXISRQTDATA[251]);
  buf B_SAXISRQTDATA252 (SAXISRQTDATA_IN[252], SAXISRQTDATA[252]);
  buf B_SAXISRQTDATA253 (SAXISRQTDATA_IN[253], SAXISRQTDATA[253]);
  buf B_SAXISRQTDATA254 (SAXISRQTDATA_IN[254], SAXISRQTDATA[254]);
  buf B_SAXISRQTDATA255 (SAXISRQTDATA_IN[255], SAXISRQTDATA[255]);
  buf B_SAXISRQTDATA26 (SAXISRQTDATA_IN[26], SAXISRQTDATA[26]);
  buf B_SAXISRQTDATA27 (SAXISRQTDATA_IN[27], SAXISRQTDATA[27]);
  buf B_SAXISRQTDATA28 (SAXISRQTDATA_IN[28], SAXISRQTDATA[28]);
  buf B_SAXISRQTDATA29 (SAXISRQTDATA_IN[29], SAXISRQTDATA[29]);
  buf B_SAXISRQTDATA3 (SAXISRQTDATA_IN[3], SAXISRQTDATA[3]);
  buf B_SAXISRQTDATA30 (SAXISRQTDATA_IN[30], SAXISRQTDATA[30]);
  buf B_SAXISRQTDATA31 (SAXISRQTDATA_IN[31], SAXISRQTDATA[31]);
  buf B_SAXISRQTDATA32 (SAXISRQTDATA_IN[32], SAXISRQTDATA[32]);
  buf B_SAXISRQTDATA33 (SAXISRQTDATA_IN[33], SAXISRQTDATA[33]);
  buf B_SAXISRQTDATA34 (SAXISRQTDATA_IN[34], SAXISRQTDATA[34]);
  buf B_SAXISRQTDATA35 (SAXISRQTDATA_IN[35], SAXISRQTDATA[35]);
  buf B_SAXISRQTDATA36 (SAXISRQTDATA_IN[36], SAXISRQTDATA[36]);
  buf B_SAXISRQTDATA37 (SAXISRQTDATA_IN[37], SAXISRQTDATA[37]);
  buf B_SAXISRQTDATA38 (SAXISRQTDATA_IN[38], SAXISRQTDATA[38]);
  buf B_SAXISRQTDATA39 (SAXISRQTDATA_IN[39], SAXISRQTDATA[39]);
  buf B_SAXISRQTDATA4 (SAXISRQTDATA_IN[4], SAXISRQTDATA[4]);
  buf B_SAXISRQTDATA40 (SAXISRQTDATA_IN[40], SAXISRQTDATA[40]);
  buf B_SAXISRQTDATA41 (SAXISRQTDATA_IN[41], SAXISRQTDATA[41]);
  buf B_SAXISRQTDATA42 (SAXISRQTDATA_IN[42], SAXISRQTDATA[42]);
  buf B_SAXISRQTDATA43 (SAXISRQTDATA_IN[43], SAXISRQTDATA[43]);
  buf B_SAXISRQTDATA44 (SAXISRQTDATA_IN[44], SAXISRQTDATA[44]);
  buf B_SAXISRQTDATA45 (SAXISRQTDATA_IN[45], SAXISRQTDATA[45]);
  buf B_SAXISRQTDATA46 (SAXISRQTDATA_IN[46], SAXISRQTDATA[46]);
  buf B_SAXISRQTDATA47 (SAXISRQTDATA_IN[47], SAXISRQTDATA[47]);
  buf B_SAXISRQTDATA48 (SAXISRQTDATA_IN[48], SAXISRQTDATA[48]);
  buf B_SAXISRQTDATA49 (SAXISRQTDATA_IN[49], SAXISRQTDATA[49]);
  buf B_SAXISRQTDATA5 (SAXISRQTDATA_IN[5], SAXISRQTDATA[5]);
  buf B_SAXISRQTDATA50 (SAXISRQTDATA_IN[50], SAXISRQTDATA[50]);
  buf B_SAXISRQTDATA51 (SAXISRQTDATA_IN[51], SAXISRQTDATA[51]);
  buf B_SAXISRQTDATA52 (SAXISRQTDATA_IN[52], SAXISRQTDATA[52]);
  buf B_SAXISRQTDATA53 (SAXISRQTDATA_IN[53], SAXISRQTDATA[53]);
  buf B_SAXISRQTDATA54 (SAXISRQTDATA_IN[54], SAXISRQTDATA[54]);
  buf B_SAXISRQTDATA55 (SAXISRQTDATA_IN[55], SAXISRQTDATA[55]);
  buf B_SAXISRQTDATA56 (SAXISRQTDATA_IN[56], SAXISRQTDATA[56]);
  buf B_SAXISRQTDATA57 (SAXISRQTDATA_IN[57], SAXISRQTDATA[57]);
  buf B_SAXISRQTDATA58 (SAXISRQTDATA_IN[58], SAXISRQTDATA[58]);
  buf B_SAXISRQTDATA59 (SAXISRQTDATA_IN[59], SAXISRQTDATA[59]);
  buf B_SAXISRQTDATA6 (SAXISRQTDATA_IN[6], SAXISRQTDATA[6]);
  buf B_SAXISRQTDATA60 (SAXISRQTDATA_IN[60], SAXISRQTDATA[60]);
  buf B_SAXISRQTDATA61 (SAXISRQTDATA_IN[61], SAXISRQTDATA[61]);
  buf B_SAXISRQTDATA62 (SAXISRQTDATA_IN[62], SAXISRQTDATA[62]);
  buf B_SAXISRQTDATA63 (SAXISRQTDATA_IN[63], SAXISRQTDATA[63]);
  buf B_SAXISRQTDATA64 (SAXISRQTDATA_IN[64], SAXISRQTDATA[64]);
  buf B_SAXISRQTDATA65 (SAXISRQTDATA_IN[65], SAXISRQTDATA[65]);
  buf B_SAXISRQTDATA66 (SAXISRQTDATA_IN[66], SAXISRQTDATA[66]);
  buf B_SAXISRQTDATA67 (SAXISRQTDATA_IN[67], SAXISRQTDATA[67]);
  buf B_SAXISRQTDATA68 (SAXISRQTDATA_IN[68], SAXISRQTDATA[68]);
  buf B_SAXISRQTDATA69 (SAXISRQTDATA_IN[69], SAXISRQTDATA[69]);
  buf B_SAXISRQTDATA7 (SAXISRQTDATA_IN[7], SAXISRQTDATA[7]);
  buf B_SAXISRQTDATA70 (SAXISRQTDATA_IN[70], SAXISRQTDATA[70]);
  buf B_SAXISRQTDATA71 (SAXISRQTDATA_IN[71], SAXISRQTDATA[71]);
  buf B_SAXISRQTDATA72 (SAXISRQTDATA_IN[72], SAXISRQTDATA[72]);
  buf B_SAXISRQTDATA73 (SAXISRQTDATA_IN[73], SAXISRQTDATA[73]);
  buf B_SAXISRQTDATA74 (SAXISRQTDATA_IN[74], SAXISRQTDATA[74]);
  buf B_SAXISRQTDATA75 (SAXISRQTDATA_IN[75], SAXISRQTDATA[75]);
  buf B_SAXISRQTDATA76 (SAXISRQTDATA_IN[76], SAXISRQTDATA[76]);
  buf B_SAXISRQTDATA77 (SAXISRQTDATA_IN[77], SAXISRQTDATA[77]);
  buf B_SAXISRQTDATA78 (SAXISRQTDATA_IN[78], SAXISRQTDATA[78]);
  buf B_SAXISRQTDATA79 (SAXISRQTDATA_IN[79], SAXISRQTDATA[79]);
  buf B_SAXISRQTDATA8 (SAXISRQTDATA_IN[8], SAXISRQTDATA[8]);
  buf B_SAXISRQTDATA80 (SAXISRQTDATA_IN[80], SAXISRQTDATA[80]);
  buf B_SAXISRQTDATA81 (SAXISRQTDATA_IN[81], SAXISRQTDATA[81]);
  buf B_SAXISRQTDATA82 (SAXISRQTDATA_IN[82], SAXISRQTDATA[82]);
  buf B_SAXISRQTDATA83 (SAXISRQTDATA_IN[83], SAXISRQTDATA[83]);
  buf B_SAXISRQTDATA84 (SAXISRQTDATA_IN[84], SAXISRQTDATA[84]);
  buf B_SAXISRQTDATA85 (SAXISRQTDATA_IN[85], SAXISRQTDATA[85]);
  buf B_SAXISRQTDATA86 (SAXISRQTDATA_IN[86], SAXISRQTDATA[86]);
  buf B_SAXISRQTDATA87 (SAXISRQTDATA_IN[87], SAXISRQTDATA[87]);
  buf B_SAXISRQTDATA88 (SAXISRQTDATA_IN[88], SAXISRQTDATA[88]);
  buf B_SAXISRQTDATA89 (SAXISRQTDATA_IN[89], SAXISRQTDATA[89]);
  buf B_SAXISRQTDATA9 (SAXISRQTDATA_IN[9], SAXISRQTDATA[9]);
  buf B_SAXISRQTDATA90 (SAXISRQTDATA_IN[90], SAXISRQTDATA[90]);
  buf B_SAXISRQTDATA91 (SAXISRQTDATA_IN[91], SAXISRQTDATA[91]);
  buf B_SAXISRQTDATA92 (SAXISRQTDATA_IN[92], SAXISRQTDATA[92]);
  buf B_SAXISRQTDATA93 (SAXISRQTDATA_IN[93], SAXISRQTDATA[93]);
  buf B_SAXISRQTDATA94 (SAXISRQTDATA_IN[94], SAXISRQTDATA[94]);
  buf B_SAXISRQTDATA95 (SAXISRQTDATA_IN[95], SAXISRQTDATA[95]);
  buf B_SAXISRQTDATA96 (SAXISRQTDATA_IN[96], SAXISRQTDATA[96]);
  buf B_SAXISRQTDATA97 (SAXISRQTDATA_IN[97], SAXISRQTDATA[97]);
  buf B_SAXISRQTDATA98 (SAXISRQTDATA_IN[98], SAXISRQTDATA[98]);
  buf B_SAXISRQTDATA99 (SAXISRQTDATA_IN[99], SAXISRQTDATA[99]);
  buf B_SAXISRQTKEEP0 (SAXISRQTKEEP_IN[0], SAXISRQTKEEP[0]);
  buf B_SAXISRQTKEEP1 (SAXISRQTKEEP_IN[1], SAXISRQTKEEP[1]);
  buf B_SAXISRQTKEEP2 (SAXISRQTKEEP_IN[2], SAXISRQTKEEP[2]);
  buf B_SAXISRQTKEEP3 (SAXISRQTKEEP_IN[3], SAXISRQTKEEP[3]);
  buf B_SAXISRQTKEEP4 (SAXISRQTKEEP_IN[4], SAXISRQTKEEP[4]);
  buf B_SAXISRQTKEEP5 (SAXISRQTKEEP_IN[5], SAXISRQTKEEP[5]);
  buf B_SAXISRQTKEEP6 (SAXISRQTKEEP_IN[6], SAXISRQTKEEP[6]);
  buf B_SAXISRQTKEEP7 (SAXISRQTKEEP_IN[7], SAXISRQTKEEP[7]);
  buf B_SAXISRQTLAST (SAXISRQTLAST_IN, SAXISRQTLAST);
  buf B_SAXISRQTUSER0 (SAXISRQTUSER_IN[0], SAXISRQTUSER[0]);
  buf B_SAXISRQTUSER1 (SAXISRQTUSER_IN[1], SAXISRQTUSER[1]);
  buf B_SAXISRQTUSER10 (SAXISRQTUSER_IN[10], SAXISRQTUSER[10]);
  buf B_SAXISRQTUSER11 (SAXISRQTUSER_IN[11], SAXISRQTUSER[11]);
  buf B_SAXISRQTUSER12 (SAXISRQTUSER_IN[12], SAXISRQTUSER[12]);
  buf B_SAXISRQTUSER13 (SAXISRQTUSER_IN[13], SAXISRQTUSER[13]);
  buf B_SAXISRQTUSER14 (SAXISRQTUSER_IN[14], SAXISRQTUSER[14]);
  buf B_SAXISRQTUSER15 (SAXISRQTUSER_IN[15], SAXISRQTUSER[15]);
  buf B_SAXISRQTUSER16 (SAXISRQTUSER_IN[16], SAXISRQTUSER[16]);
  buf B_SAXISRQTUSER17 (SAXISRQTUSER_IN[17], SAXISRQTUSER[17]);
  buf B_SAXISRQTUSER18 (SAXISRQTUSER_IN[18], SAXISRQTUSER[18]);
  buf B_SAXISRQTUSER19 (SAXISRQTUSER_IN[19], SAXISRQTUSER[19]);
  buf B_SAXISRQTUSER2 (SAXISRQTUSER_IN[2], SAXISRQTUSER[2]);
  buf B_SAXISRQTUSER20 (SAXISRQTUSER_IN[20], SAXISRQTUSER[20]);
  buf B_SAXISRQTUSER21 (SAXISRQTUSER_IN[21], SAXISRQTUSER[21]);
  buf B_SAXISRQTUSER22 (SAXISRQTUSER_IN[22], SAXISRQTUSER[22]);
  buf B_SAXISRQTUSER23 (SAXISRQTUSER_IN[23], SAXISRQTUSER[23]);
  buf B_SAXISRQTUSER24 (SAXISRQTUSER_IN[24], SAXISRQTUSER[24]);
  buf B_SAXISRQTUSER25 (SAXISRQTUSER_IN[25], SAXISRQTUSER[25]);
  buf B_SAXISRQTUSER26 (SAXISRQTUSER_IN[26], SAXISRQTUSER[26]);
  buf B_SAXISRQTUSER27 (SAXISRQTUSER_IN[27], SAXISRQTUSER[27]);
  buf B_SAXISRQTUSER28 (SAXISRQTUSER_IN[28], SAXISRQTUSER[28]);
  buf B_SAXISRQTUSER29 (SAXISRQTUSER_IN[29], SAXISRQTUSER[29]);
  buf B_SAXISRQTUSER3 (SAXISRQTUSER_IN[3], SAXISRQTUSER[3]);
  buf B_SAXISRQTUSER30 (SAXISRQTUSER_IN[30], SAXISRQTUSER[30]);
  buf B_SAXISRQTUSER31 (SAXISRQTUSER_IN[31], SAXISRQTUSER[31]);
  buf B_SAXISRQTUSER32 (SAXISRQTUSER_IN[32], SAXISRQTUSER[32]);
  buf B_SAXISRQTUSER33 (SAXISRQTUSER_IN[33], SAXISRQTUSER[33]);
  buf B_SAXISRQTUSER34 (SAXISRQTUSER_IN[34], SAXISRQTUSER[34]);
  buf B_SAXISRQTUSER35 (SAXISRQTUSER_IN[35], SAXISRQTUSER[35]);
  buf B_SAXISRQTUSER36 (SAXISRQTUSER_IN[36], SAXISRQTUSER[36]);
  buf B_SAXISRQTUSER37 (SAXISRQTUSER_IN[37], SAXISRQTUSER[37]);
  buf B_SAXISRQTUSER38 (SAXISRQTUSER_IN[38], SAXISRQTUSER[38]);
  buf B_SAXISRQTUSER39 (SAXISRQTUSER_IN[39], SAXISRQTUSER[39]);
  buf B_SAXISRQTUSER4 (SAXISRQTUSER_IN[4], SAXISRQTUSER[4]);
  buf B_SAXISRQTUSER40 (SAXISRQTUSER_IN[40], SAXISRQTUSER[40]);
  buf B_SAXISRQTUSER41 (SAXISRQTUSER_IN[41], SAXISRQTUSER[41]);
  buf B_SAXISRQTUSER42 (SAXISRQTUSER_IN[42], SAXISRQTUSER[42]);
  buf B_SAXISRQTUSER43 (SAXISRQTUSER_IN[43], SAXISRQTUSER[43]);
  buf B_SAXISRQTUSER44 (SAXISRQTUSER_IN[44], SAXISRQTUSER[44]);
  buf B_SAXISRQTUSER45 (SAXISRQTUSER_IN[45], SAXISRQTUSER[45]);
  buf B_SAXISRQTUSER46 (SAXISRQTUSER_IN[46], SAXISRQTUSER[46]);
  buf B_SAXISRQTUSER47 (SAXISRQTUSER_IN[47], SAXISRQTUSER[47]);
  buf B_SAXISRQTUSER48 (SAXISRQTUSER_IN[48], SAXISRQTUSER[48]);
  buf B_SAXISRQTUSER49 (SAXISRQTUSER_IN[49], SAXISRQTUSER[49]);
  buf B_SAXISRQTUSER5 (SAXISRQTUSER_IN[5], SAXISRQTUSER[5]);
  buf B_SAXISRQTUSER50 (SAXISRQTUSER_IN[50], SAXISRQTUSER[50]);
  buf B_SAXISRQTUSER51 (SAXISRQTUSER_IN[51], SAXISRQTUSER[51]);
  buf B_SAXISRQTUSER52 (SAXISRQTUSER_IN[52], SAXISRQTUSER[52]);
  buf B_SAXISRQTUSER53 (SAXISRQTUSER_IN[53], SAXISRQTUSER[53]);
  buf B_SAXISRQTUSER54 (SAXISRQTUSER_IN[54], SAXISRQTUSER[54]);
  buf B_SAXISRQTUSER55 (SAXISRQTUSER_IN[55], SAXISRQTUSER[55]);
  buf B_SAXISRQTUSER56 (SAXISRQTUSER_IN[56], SAXISRQTUSER[56]);
  buf B_SAXISRQTUSER57 (SAXISRQTUSER_IN[57], SAXISRQTUSER[57]);
  buf B_SAXISRQTUSER58 (SAXISRQTUSER_IN[58], SAXISRQTUSER[58]);
  buf B_SAXISRQTUSER59 (SAXISRQTUSER_IN[59], SAXISRQTUSER[59]);
  buf B_SAXISRQTUSER6 (SAXISRQTUSER_IN[6], SAXISRQTUSER[6]);
  buf B_SAXISRQTUSER7 (SAXISRQTUSER_IN[7], SAXISRQTUSER[7]);
  buf B_SAXISRQTUSER8 (SAXISRQTUSER_IN[8], SAXISRQTUSER[8]);
  buf B_SAXISRQTUSER9 (SAXISRQTUSER_IN[9], SAXISRQTUSER[9]);
  buf B_SAXISRQTVALID (SAXISRQTVALID_IN, SAXISRQTVALID);
  buf B_USERCLK (USERCLK_IN, USERCLK);

  wire [11:0] delay_CFGFCCPLD;
  wire [11:0] delay_CFGFCNPD;
  wire [11:0] delay_CFGFCPD;
  wire [11:0] delay_CFGVFSTATUS;
  wire [143:0] delay_MIREPLAYRAMWRITEDATA;
  wire [143:0] delay_MIREQUESTRAMWRITEDATA;
  wire [15:0] delay_CFGPERFUNCSTATUSDATA;
  wire [15:0] delay_DBGDATAOUT;
  wire [15:0] delay_DRPDO;
  wire [17:0] delay_CFGVFPOWERSTATE;
  wire [17:0] delay_CFGVFTPHSTMODE;
  wire [1:0] delay_CFGDPASUBSTATECHANGE;
  wire [1:0] delay_CFGFLRINPROCESS;
  wire [1:0] delay_CFGINTERRUPTMSIENABLE;
  wire [1:0] delay_CFGINTERRUPTMSIXENABLE;
  wire [1:0] delay_CFGINTERRUPTMSIXMASK;
  wire [1:0] delay_CFGLINKPOWERSTATE;
  wire [1:0] delay_CFGOBFFENABLE;
  wire [1:0] delay_CFGPHYLINKSTATUS;
  wire [1:0] delay_CFGRCBSTATUS;
  wire [1:0] delay_CFGTPHREQUESTERENABLE;
  wire [1:0] delay_MIREPLAYRAMREADENABLE;
  wire [1:0] delay_MIREPLAYRAMWRITEENABLE;
  wire [1:0] delay_PCIERQTAGAV;
  wire [1:0] delay_PCIETFCNPDAV;
  wire [1:0] delay_PCIETFCNPHAV;
  wire [1:0] delay_PIPERX0EQCONTROL;
  wire [1:0] delay_PIPERX1EQCONTROL;
  wire [1:0] delay_PIPERX2EQCONTROL;
  wire [1:0] delay_PIPERX3EQCONTROL;
  wire [1:0] delay_PIPERX4EQCONTROL;
  wire [1:0] delay_PIPERX5EQCONTROL;
  wire [1:0] delay_PIPERX6EQCONTROL;
  wire [1:0] delay_PIPERX7EQCONTROL;
  wire [1:0] delay_PIPETX0CHARISK;
  wire [1:0] delay_PIPETX0EQCONTROL;
  wire [1:0] delay_PIPETX0POWERDOWN;
  wire [1:0] delay_PIPETX0SYNCHEADER;
  wire [1:0] delay_PIPETX1CHARISK;
  wire [1:0] delay_PIPETX1EQCONTROL;
  wire [1:0] delay_PIPETX1POWERDOWN;
  wire [1:0] delay_PIPETX1SYNCHEADER;
  wire [1:0] delay_PIPETX2CHARISK;
  wire [1:0] delay_PIPETX2EQCONTROL;
  wire [1:0] delay_PIPETX2POWERDOWN;
  wire [1:0] delay_PIPETX2SYNCHEADER;
  wire [1:0] delay_PIPETX3CHARISK;
  wire [1:0] delay_PIPETX3EQCONTROL;
  wire [1:0] delay_PIPETX3POWERDOWN;
  wire [1:0] delay_PIPETX3SYNCHEADER;
  wire [1:0] delay_PIPETX4CHARISK;
  wire [1:0] delay_PIPETX4EQCONTROL;
  wire [1:0] delay_PIPETX4POWERDOWN;
  wire [1:0] delay_PIPETX4SYNCHEADER;
  wire [1:0] delay_PIPETX5CHARISK;
  wire [1:0] delay_PIPETX5EQCONTROL;
  wire [1:0] delay_PIPETX5POWERDOWN;
  wire [1:0] delay_PIPETX5SYNCHEADER;
  wire [1:0] delay_PIPETX6CHARISK;
  wire [1:0] delay_PIPETX6EQCONTROL;
  wire [1:0] delay_PIPETX6POWERDOWN;
  wire [1:0] delay_PIPETX6SYNCHEADER;
  wire [1:0] delay_PIPETX7CHARISK;
  wire [1:0] delay_PIPETX7EQCONTROL;
  wire [1:0] delay_PIPETX7POWERDOWN;
  wire [1:0] delay_PIPETX7SYNCHEADER;
  wire [1:0] delay_PIPETXRATE;
  wire [1:0] delay_PLEQPHASE;
  wire [255:0] delay_MAXISCQTDATA;
  wire [255:0] delay_MAXISRCTDATA;
  wire [2:0] delay_CFGCURRENTSPEED;
  wire [2:0] delay_CFGMAXPAYLOAD;
  wire [2:0] delay_CFGMAXREADREQ;
  wire [2:0] delay_CFGTPHFUNCTIONNUM;
  wire [2:0] delay_PIPERX0EQPRESET;
  wire [2:0] delay_PIPERX1EQPRESET;
  wire [2:0] delay_PIPERX2EQPRESET;
  wire [2:0] delay_PIPERX3EQPRESET;
  wire [2:0] delay_PIPERX4EQPRESET;
  wire [2:0] delay_PIPERX5EQPRESET;
  wire [2:0] delay_PIPERX6EQPRESET;
  wire [2:0] delay_PIPERX7EQPRESET;
  wire [2:0] delay_PIPETXMARGIN;
  wire [31:0] delay_CFGEXTWRITEDATA;
  wire [31:0] delay_CFGINTERRUPTMSIDATA;
  wire [31:0] delay_CFGMGMTREADDATA;
  wire [31:0] delay_CFGTPHSTTWRITEDATA;
  wire [31:0] delay_PIPETX0DATA;
  wire [31:0] delay_PIPETX1DATA;
  wire [31:0] delay_PIPETX2DATA;
  wire [31:0] delay_PIPETX3DATA;
  wire [31:0] delay_PIPETX4DATA;
  wire [31:0] delay_PIPETX5DATA;
  wire [31:0] delay_PIPETX6DATA;
  wire [31:0] delay_PIPETX7DATA;
  wire [3:0] delay_CFGEXTWRITEBYTEENABLE;
  wire [3:0] delay_CFGNEGOTIATEDWIDTH;
  wire [3:0] delay_CFGTPHSTTWRITEBYTEVALID;
  wire [3:0] delay_MICOMPLETIONRAMREADENABLEL;
  wire [3:0] delay_MICOMPLETIONRAMREADENABLEU;
  wire [3:0] delay_MICOMPLETIONRAMWRITEENABLEL;
  wire [3:0] delay_MICOMPLETIONRAMWRITEENABLEU;
  wire [3:0] delay_MIREQUESTRAMREADENABLE;
  wire [3:0] delay_MIREQUESTRAMWRITEENABLE;
  wire [3:0] delay_PCIERQSEQNUM;
  wire [3:0] delay_PIPERX0EQLPTXPRESET;
  wire [3:0] delay_PIPERX1EQLPTXPRESET;
  wire [3:0] delay_PIPERX2EQLPTXPRESET;
  wire [3:0] delay_PIPERX3EQLPTXPRESET;
  wire [3:0] delay_PIPERX4EQLPTXPRESET;
  wire [3:0] delay_PIPERX5EQLPTXPRESET;
  wire [3:0] delay_PIPERX6EQLPTXPRESET;
  wire [3:0] delay_PIPERX7EQLPTXPRESET;
  wire [3:0] delay_PIPETX0EQPRESET;
  wire [3:0] delay_PIPETX1EQPRESET;
  wire [3:0] delay_PIPETX2EQPRESET;
  wire [3:0] delay_PIPETX3EQPRESET;
  wire [3:0] delay_PIPETX4EQPRESET;
  wire [3:0] delay_PIPETX5EQPRESET;
  wire [3:0] delay_PIPETX6EQPRESET;
  wire [3:0] delay_PIPETX7EQPRESET;
  wire [3:0] delay_SAXISCCTREADY;
  wire [3:0] delay_SAXISRQTREADY;
  wire [4:0] delay_CFGMSGRECEIVEDTYPE;
  wire [4:0] delay_CFGTPHSTTADDRESS;
  wire [5:0] delay_CFGFUNCTIONPOWERSTATE;
  wire [5:0] delay_CFGINTERRUPTMSIMMENABLE;
  wire [5:0] delay_CFGINTERRUPTMSIVFENABLE;
  wire [5:0] delay_CFGINTERRUPTMSIXVFENABLE;
  wire [5:0] delay_CFGINTERRUPTMSIXVFMASK;
  wire [5:0] delay_CFGLTSSMSTATE;
  wire [5:0] delay_CFGTPHSTMODE;
  wire [5:0] delay_CFGVFFLRINPROCESS;
  wire [5:0] delay_CFGVFTPHREQUESTERENABLE;
  wire [5:0] delay_PCIECQNPREQCOUNT;
  wire [5:0] delay_PCIERQTAG;
  wire [5:0] delay_PIPERX0EQLPLFFS;
  wire [5:0] delay_PIPERX1EQLPLFFS;
  wire [5:0] delay_PIPERX2EQLPLFFS;
  wire [5:0] delay_PIPERX3EQLPLFFS;
  wire [5:0] delay_PIPERX4EQLPLFFS;
  wire [5:0] delay_PIPERX5EQLPLFFS;
  wire [5:0] delay_PIPERX6EQLPLFFS;
  wire [5:0] delay_PIPERX7EQLPLFFS;
  wire [5:0] delay_PIPETX0EQDEEMPH;
  wire [5:0] delay_PIPETX1EQDEEMPH;
  wire [5:0] delay_PIPETX2EQDEEMPH;
  wire [5:0] delay_PIPETX3EQDEEMPH;
  wire [5:0] delay_PIPETX4EQDEEMPH;
  wire [5:0] delay_PIPETX5EQDEEMPH;
  wire [5:0] delay_PIPETX6EQDEEMPH;
  wire [5:0] delay_PIPETX7EQDEEMPH;
  wire [71:0] delay_MICOMPLETIONRAMWRITEDATAL;
  wire [71:0] delay_MICOMPLETIONRAMWRITEDATAU;
  wire [74:0] delay_MAXISRCTUSER;
  wire [7:0] delay_CFGEXTFUNCTIONNUMBER;
  wire [7:0] delay_CFGFCCPLH;
  wire [7:0] delay_CFGFCNPH;
  wire [7:0] delay_CFGFCPH;
  wire [7:0] delay_CFGFUNCTIONSTATUS;
  wire [7:0] delay_CFGMSGRECEIVEDDATA;
  wire [7:0] delay_MAXISCQTKEEP;
  wire [7:0] delay_MAXISRCTKEEP;
  wire [7:0] delay_PLGEN3PCSRXSLIDE;
  wire [84:0] delay_MAXISCQTUSER;
  wire [8:0] delay_MIREPLAYRAMADDRESS;
  wire [8:0] delay_MIREQUESTRAMREADADDRESSA;
  wire [8:0] delay_MIREQUESTRAMREADADDRESSB;
  wire [8:0] delay_MIREQUESTRAMWRITEADDRESSA;
  wire [8:0] delay_MIREQUESTRAMWRITEADDRESSB;
  wire [9:0] delay_CFGEXTREGISTERNUMBER;
  wire [9:0] delay_MICOMPLETIONRAMREADADDRESSAL;
  wire [9:0] delay_MICOMPLETIONRAMREADADDRESSAU;
  wire [9:0] delay_MICOMPLETIONRAMREADADDRESSBL;
  wire [9:0] delay_MICOMPLETIONRAMREADADDRESSBU;
  wire [9:0] delay_MICOMPLETIONRAMWRITEADDRESSAL;
  wire [9:0] delay_MICOMPLETIONRAMWRITEADDRESSAU;
  wire [9:0] delay_MICOMPLETIONRAMWRITEADDRESSBL;
  wire [9:0] delay_MICOMPLETIONRAMWRITEADDRESSBU;
  wire delay_CFGERRCOROUT;
  wire delay_CFGERRFATALOUT;
  wire delay_CFGERRNONFATALOUT;
  wire delay_CFGEXTREADRECEIVED;
  wire delay_CFGEXTWRITERECEIVED;
  wire delay_CFGHOTRESETOUT;
  wire delay_CFGINPUTUPDATEDONE;
  wire delay_CFGINTERRUPTAOUTPUT;
  wire delay_CFGINTERRUPTBOUTPUT;
  wire delay_CFGINTERRUPTCOUTPUT;
  wire delay_CFGINTERRUPTDOUTPUT;
  wire delay_CFGINTERRUPTMSIFAIL;
  wire delay_CFGINTERRUPTMSIMASKUPDATE;
  wire delay_CFGINTERRUPTMSISENT;
  wire delay_CFGINTERRUPTMSIXFAIL;
  wire delay_CFGINTERRUPTMSIXSENT;
  wire delay_CFGINTERRUPTSENT;
  wire delay_CFGLOCALERROR;
  wire delay_CFGLTRENABLE;
  wire delay_CFGMCUPDATEDONE;
  wire delay_CFGMGMTREADWRITEDONE;
  wire delay_CFGMSGRECEIVED;
  wire delay_CFGMSGTRANSMITDONE;
  wire delay_CFGPERFUNCTIONUPDATEDONE;
  wire delay_CFGPHYLINKDOWN;
  wire delay_CFGPLSTATUSCHANGE;
  wire delay_CFGPOWERSTATECHANGEINTERRUPT;
  wire delay_CFGTPHSTTREADENABLE;
  wire delay_CFGTPHSTTWRITEENABLE;
  wire delay_DRPRDY;
  wire delay_MAXISCQTLAST;
  wire delay_MAXISCQTVALID;
  wire delay_MAXISRCTLAST;
  wire delay_MAXISRCTVALID;
  wire delay_PCIERQSEQNUMVLD;
  wire delay_PCIERQTAGVLD;
  wire delay_PIPERX0POLARITY;
  wire delay_PIPERX1POLARITY;
  wire delay_PIPERX2POLARITY;
  wire delay_PIPERX3POLARITY;
  wire delay_PIPERX4POLARITY;
  wire delay_PIPERX5POLARITY;
  wire delay_PIPERX6POLARITY;
  wire delay_PIPERX7POLARITY;
  wire delay_PIPETX0COMPLIANCE;
  wire delay_PIPETX0DATAVALID;
  wire delay_PIPETX0ELECIDLE;
  wire delay_PIPETX0STARTBLOCK;
  wire delay_PIPETX1COMPLIANCE;
  wire delay_PIPETX1DATAVALID;
  wire delay_PIPETX1ELECIDLE;
  wire delay_PIPETX1STARTBLOCK;
  wire delay_PIPETX2COMPLIANCE;
  wire delay_PIPETX2DATAVALID;
  wire delay_PIPETX2ELECIDLE;
  wire delay_PIPETX2STARTBLOCK;
  wire delay_PIPETX3COMPLIANCE;
  wire delay_PIPETX3DATAVALID;
  wire delay_PIPETX3ELECIDLE;
  wire delay_PIPETX3STARTBLOCK;
  wire delay_PIPETX4COMPLIANCE;
  wire delay_PIPETX4DATAVALID;
  wire delay_PIPETX4ELECIDLE;
  wire delay_PIPETX4STARTBLOCK;
  wire delay_PIPETX5COMPLIANCE;
  wire delay_PIPETX5DATAVALID;
  wire delay_PIPETX5ELECIDLE;
  wire delay_PIPETX5STARTBLOCK;
  wire delay_PIPETX6COMPLIANCE;
  wire delay_PIPETX6DATAVALID;
  wire delay_PIPETX6ELECIDLE;
  wire delay_PIPETX6STARTBLOCK;
  wire delay_PIPETX7COMPLIANCE;
  wire delay_PIPETX7DATAVALID;
  wire delay_PIPETX7ELECIDLE;
  wire delay_PIPETX7STARTBLOCK;
  wire delay_PIPETXDEEMPH;
  wire delay_PIPETXRCVRDET;
  wire delay_PIPETXRESET;
  wire delay_PIPETXSWING;
  wire delay_PLEQINPROGRESS;

  wire [10:0] delay_DRPADDR;
  wire [143:0] delay_MICOMPLETIONRAMREADDATA;
  wire [143:0] delay_MIREPLAYRAMREADDATA;
  wire [143:0] delay_MIREQUESTRAMREADDATA;
  wire [15:0] delay_CFGDEVID;
  wire [15:0] delay_CFGSUBSYSID;
  wire [15:0] delay_CFGSUBSYSVENDID;
  wire [15:0] delay_CFGVENDID;
  wire [15:0] delay_DRPDI;
  wire [17:0] delay_PIPERX0EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX1EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX2EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX3EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX4EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX5EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX6EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPERX7EQLPNEWTXCOEFFORPRESET;
  wire [17:0] delay_PIPETX0EQCOEFF;
  wire [17:0] delay_PIPETX1EQCOEFF;
  wire [17:0] delay_PIPETX2EQCOEFF;
  wire [17:0] delay_PIPETX3EQCOEFF;
  wire [17:0] delay_PIPETX4EQCOEFF;
  wire [17:0] delay_PIPETX5EQCOEFF;
  wire [17:0] delay_PIPETX6EQCOEFF;
  wire [17:0] delay_PIPETX7EQCOEFF;
  wire [18:0] delay_CFGMGMTADDR;
  wire [1:0] delay_CFGFLRDONE;
  wire [1:0] delay_CFGINTERRUPTMSITPHTYPE;
  wire [1:0] delay_CFGINTERRUPTPENDING;
  wire [1:0] delay_PIPERX0CHARISK;
  wire [1:0] delay_PIPERX0SYNCHEADER;
  wire [1:0] delay_PIPERX1CHARISK;
  wire [1:0] delay_PIPERX1SYNCHEADER;
  wire [1:0] delay_PIPERX2CHARISK;
  wire [1:0] delay_PIPERX2SYNCHEADER;
  wire [1:0] delay_PIPERX3CHARISK;
  wire [1:0] delay_PIPERX3SYNCHEADER;
  wire [1:0] delay_PIPERX4CHARISK;
  wire [1:0] delay_PIPERX4SYNCHEADER;
  wire [1:0] delay_PIPERX5CHARISK;
  wire [1:0] delay_PIPERX5SYNCHEADER;
  wire [1:0] delay_PIPERX6CHARISK;
  wire [1:0] delay_PIPERX6SYNCHEADER;
  wire [1:0] delay_PIPERX7CHARISK;
  wire [1:0] delay_PIPERX7SYNCHEADER;
  wire [21:0] delay_MAXISCQTREADY;
  wire [21:0] delay_MAXISRCTREADY;
  wire [255:0] delay_SAXISCCTDATA;
  wire [255:0] delay_SAXISRQTDATA;
  wire [2:0] delay_CFGDSFUNCTIONNUMBER;
  wire [2:0] delay_CFGFCSEL;
  wire [2:0] delay_CFGINTERRUPTMSIATTR;
  wire [2:0] delay_CFGINTERRUPTMSIFUNCTIONNUMBER;
  wire [2:0] delay_CFGMSGTRANSMITTYPE;
  wire [2:0] delay_CFGPERFUNCSTATUSCONTROL;
  wire [2:0] delay_CFGPERFUNCTIONNUMBER;
  wire [2:0] delay_PIPERX0STATUS;
  wire [2:0] delay_PIPERX1STATUS;
  wire [2:0] delay_PIPERX2STATUS;
  wire [2:0] delay_PIPERX3STATUS;
  wire [2:0] delay_PIPERX4STATUS;
  wire [2:0] delay_PIPERX5STATUS;
  wire [2:0] delay_PIPERX6STATUS;
  wire [2:0] delay_PIPERX7STATUS;
  wire [31:0] delay_CFGEXTREADDATA;
  wire [31:0] delay_CFGINTERRUPTMSIINT;
  wire [31:0] delay_CFGINTERRUPTMSIXDATA;
  wire [31:0] delay_CFGMGMTWRITEDATA;
  wire [31:0] delay_CFGMSGTRANSMITDATA;
  wire [31:0] delay_CFGTPHSTTREADDATA;
  wire [31:0] delay_PIPERX0DATA;
  wire [31:0] delay_PIPERX1DATA;
  wire [31:0] delay_PIPERX2DATA;
  wire [31:0] delay_PIPERX3DATA;
  wire [31:0] delay_PIPERX4DATA;
  wire [31:0] delay_PIPERX5DATA;
  wire [31:0] delay_PIPERX6DATA;
  wire [31:0] delay_PIPERX7DATA;
  wire [32:0] delay_SAXISCCTUSER;
  wire [3:0] delay_CFGINTERRUPTINT;
  wire [3:0] delay_CFGINTERRUPTMSISELECT;
  wire [3:0] delay_CFGMGMTBYTEENABLE;
  wire [4:0] delay_CFGDSDEVICENUMBER;
  wire [59:0] delay_SAXISRQTUSER;
  wire [5:0] delay_CFGVFFLRDONE;
  wire [5:0] delay_PIPEEQFS;
  wire [5:0] delay_PIPEEQLF;
  wire [63:0] delay_CFGDSN;
  wire [63:0] delay_CFGINTERRUPTMSIPENDINGSTATUS;
  wire [63:0] delay_CFGINTERRUPTMSIXADDRESS;
  wire [7:0] delay_CFGDSBUSNUMBER;
  wire [7:0] delay_CFGDSPORTNUMBER;
  wire [7:0] delay_CFGREVID;
  wire [7:0] delay_PLGEN3PCSRXSYNCDONE;
  wire [7:0] delay_SAXISCCTKEEP;
  wire [7:0] delay_SAXISRQTKEEP;
  wire [8:0] delay_CFGINTERRUPTMSITPHSTTAG;
  wire delay_CFGCONFIGSPACEENABLE;
  wire delay_CFGERRCORIN;
  wire delay_CFGERRUNCORIN;
  wire delay_CFGEXTREADDATAVALID;
  wire delay_CFGHOTRESETIN;
  wire delay_CFGINPUTUPDATEREQUEST;
  wire delay_CFGINTERRUPTMSITPHPRESENT;
  wire delay_CFGINTERRUPTMSIXINT;
  wire delay_CFGLINKTRAININGENABLE;
  wire delay_CFGMCUPDATEREQUEST;
  wire delay_CFGMGMTREAD;
  wire delay_CFGMGMTTYPE1CFGREGACCESS;
  wire delay_CFGMGMTWRITE;
  wire delay_CFGMSGTRANSMIT;
  wire delay_CFGPERFUNCTIONOUTPUTREQUEST;
  wire delay_CFGPOWERSTATECHANGEACK;
  wire delay_CFGREQPMTRANSITIONL23READY;
  wire delay_CFGTPHSTTREADDATAVALID;
  wire delay_CORECLK;
  wire delay_CORECLKMICOMPLETIONRAML;
  wire delay_CORECLKMICOMPLETIONRAMU;
  wire delay_CORECLKMIREPLAYRAM;
  wire delay_CORECLKMIREQUESTRAM;
  wire delay_DRPCLK;
  wire delay_DRPEN;
  wire delay_DRPWE;
  wire delay_MGMTRESETN;
  wire delay_MGMTSTICKYRESETN;
  wire delay_PCIECQNPREQ;
  wire delay_PIPECLK;
  wire delay_PIPERESETN;
  wire delay_PIPERX0DATAVALID;
  wire delay_PIPERX0ELECIDLE;
  wire delay_PIPERX0EQDONE;
  wire delay_PIPERX0EQLPADAPTDONE;
  wire delay_PIPERX0EQLPLFFSSEL;
  wire delay_PIPERX0PHYSTATUS;
  wire delay_PIPERX0STARTBLOCK;
  wire delay_PIPERX0VALID;
  wire delay_PIPERX1DATAVALID;
  wire delay_PIPERX1ELECIDLE;
  wire delay_PIPERX1EQDONE;
  wire delay_PIPERX1EQLPADAPTDONE;
  wire delay_PIPERX1EQLPLFFSSEL;
  wire delay_PIPERX1PHYSTATUS;
  wire delay_PIPERX1STARTBLOCK;
  wire delay_PIPERX1VALID;
  wire delay_PIPERX2DATAVALID;
  wire delay_PIPERX2ELECIDLE;
  wire delay_PIPERX2EQDONE;
  wire delay_PIPERX2EQLPADAPTDONE;
  wire delay_PIPERX2EQLPLFFSSEL;
  wire delay_PIPERX2PHYSTATUS;
  wire delay_PIPERX2STARTBLOCK;
  wire delay_PIPERX2VALID;
  wire delay_PIPERX3DATAVALID;
  wire delay_PIPERX3ELECIDLE;
  wire delay_PIPERX3EQDONE;
  wire delay_PIPERX3EQLPADAPTDONE;
  wire delay_PIPERX3EQLPLFFSSEL;
  wire delay_PIPERX3PHYSTATUS;
  wire delay_PIPERX3STARTBLOCK;
  wire delay_PIPERX3VALID;
  wire delay_PIPERX4DATAVALID;
  wire delay_PIPERX4ELECIDLE;
  wire delay_PIPERX4EQDONE;
  wire delay_PIPERX4EQLPADAPTDONE;
  wire delay_PIPERX4EQLPLFFSSEL;
  wire delay_PIPERX4PHYSTATUS;
  wire delay_PIPERX4STARTBLOCK;
  wire delay_PIPERX4VALID;
  wire delay_PIPERX5DATAVALID;
  wire delay_PIPERX5ELECIDLE;
  wire delay_PIPERX5EQDONE;
  wire delay_PIPERX5EQLPADAPTDONE;
  wire delay_PIPERX5EQLPLFFSSEL;
  wire delay_PIPERX5PHYSTATUS;
  wire delay_PIPERX5STARTBLOCK;
  wire delay_PIPERX5VALID;
  wire delay_PIPERX6DATAVALID;
  wire delay_PIPERX6ELECIDLE;
  wire delay_PIPERX6EQDONE;
  wire delay_PIPERX6EQLPADAPTDONE;
  wire delay_PIPERX6EQLPLFFSSEL;
  wire delay_PIPERX6PHYSTATUS;
  wire delay_PIPERX6STARTBLOCK;
  wire delay_PIPERX6VALID;
  wire delay_PIPERX7DATAVALID;
  wire delay_PIPERX7ELECIDLE;
  wire delay_PIPERX7EQDONE;
  wire delay_PIPERX7EQLPADAPTDONE;
  wire delay_PIPERX7EQLPLFFSSEL;
  wire delay_PIPERX7PHYSTATUS;
  wire delay_PIPERX7STARTBLOCK;
  wire delay_PIPERX7VALID;
  wire delay_PIPETX0EQDONE;
  wire delay_PIPETX1EQDONE;
  wire delay_PIPETX2EQDONE;
  wire delay_PIPETX3EQDONE;
  wire delay_PIPETX4EQDONE;
  wire delay_PIPETX5EQDONE;
  wire delay_PIPETX6EQDONE;
  wire delay_PIPETX7EQDONE;
  wire delay_PLDISABLESCRAMBLER;
  wire delay_PLEQRESETEIEOSCOUNT;
  wire delay_PLGEN3PCSDISABLE;
  wire delay_RECCLK;
  wire delay_RESETN;
  wire delay_SAXISCCTLAST;
  wire delay_SAXISCCTVALID;
  wire delay_SAXISRQTLAST;
  wire delay_SAXISRQTVALID;
  wire delay_USERCLK;


   //drp monitor
   reg drpen_r1 = 1'b0;
   reg drpen_r2 = 1'b0;
   reg drpwe_r1 = 1'b0;
   reg drpwe_r2 = 1'b0;
   
   reg [1:0] sfsm = 2'b01;
    
   localparam FSM_IDLE = 2'b01;  
   localparam FSM_WAIT = 2'b10;
  

   always @(posedge delay_DRPCLK)
     begin
	// pipeline the DRPEN and DRPWE
        drpen_r1 <= delay_DRPEN;
        drpwe_r1 <= delay_DRPWE;
	drpen_r2 <= drpen_r1;
        drpwe_r2 <= drpwe_r1;

	
	// Check -  if DRPEN or DRPWE is more than 1 DCLK
	if ((drpen_r1 == 1'b1) && (drpen_r2 == 1'b1)) 
	  begin
	     $display("DRC Error : DRPEN is high for more than 1 DRPCLK on %m instance");
	     $finish; 
          end
	
	if ((drpwe_r1 == 1'b1) && (drpwe_r2 == 1'b1))
	  begin
             $display("DRC Error : DRPWE is high for more than 1 DRPCLK on %m instance");
             $finish;
          end


	//After the 1st DRPEN pulse, check the DRPEN and DRPRDY.
	case (sfsm)
          FSM_IDLE:   
            begin
               if(delay_DRPEN == 1'b1)
		 sfsm <= FSM_WAIT;  
            end
          
          FSM_WAIT:
            begin
               // After the 1st DRPEN, 4 cases can happen
               // DRPEN DRPRDY NEXT STATE
               // 0     0      FSM_WAIT - wait for DRPRDY
               // 0     1      FSM_IDLE - normal operation
               // 1     0      FSM_WAIT - display error and wait for DRPRDY
               // 1     1      FSM_WAIT - normal operation. Per UG470, DRPEN and DRPRDY can be at the same cycle.
               
               //Add the check for another DPREN pulse
               if(delay_DRPEN === 1'b1 && delay_DRPRDY === 1'b0) 
		 begin
		    $display("DRC Error : DRPEN is enabled before DRPRDY returns on %m instance");  
		    $finish;
		 end

               //Add the check for another DRPWE pulse
               if ((delay_DRPWE === 1'b1) && (delay_DRPEN === 1'b0))
		 begin
		    $display("DRC Error : DRPWE is enabled before DRPRDY returns on %m instance");
		    $finish;
		 end
                    
               if ((delay_DRPRDY === 1'b1) && (delay_DRPEN === 1'b0))
		 begin
		    sfsm <= FSM_IDLE;
		 end  
               
               if ((delay_DRPRDY === 1'b1)&& (delay_DRPEN === 1'b1))
		 begin
		    sfsm <= FSM_WAIT;
		 end  
            end
        
          default:                  
            begin
               $display("DRC Error : Default state in DRP FSM.");
               $finish;
            end
	endcase

     end // always @ (posedge delay_DRPCLK)
   //end drp monitor      

   
  assign #(out_delay) CFGCURRENTSPEED_OUT = delay_CFGCURRENTSPEED;
  assign #(out_delay) CFGDPASUBSTATECHANGE_OUT = delay_CFGDPASUBSTATECHANGE;
  assign #(out_delay) CFGERRCOROUT_OUT = delay_CFGERRCOROUT;
  assign #(out_delay) CFGERRFATALOUT_OUT = delay_CFGERRFATALOUT;
  assign #(out_delay) CFGERRNONFATALOUT_OUT = delay_CFGERRNONFATALOUT;
  assign #(out_delay) CFGEXTFUNCTIONNUMBER_OUT = delay_CFGEXTFUNCTIONNUMBER;
  assign #(out_delay) CFGEXTREADRECEIVED_OUT = delay_CFGEXTREADRECEIVED;
  assign #(out_delay) CFGEXTREGISTERNUMBER_OUT = delay_CFGEXTREGISTERNUMBER;
  assign #(out_delay) CFGEXTWRITEBYTEENABLE_OUT = delay_CFGEXTWRITEBYTEENABLE;
  assign #(out_delay) CFGEXTWRITEDATA_OUT = delay_CFGEXTWRITEDATA;
  assign #(out_delay) CFGEXTWRITERECEIVED_OUT = delay_CFGEXTWRITERECEIVED;
  assign #(out_delay) CFGFCCPLD_OUT = delay_CFGFCCPLD;
  assign #(out_delay) CFGFCCPLH_OUT = delay_CFGFCCPLH;
  assign #(out_delay) CFGFCNPD_OUT = delay_CFGFCNPD;
  assign #(out_delay) CFGFCNPH_OUT = delay_CFGFCNPH;
  assign #(out_delay) CFGFCPD_OUT = delay_CFGFCPD;
  assign #(out_delay) CFGFCPH_OUT = delay_CFGFCPH;
  assign #(out_delay) CFGFLRINPROCESS_OUT = delay_CFGFLRINPROCESS;
  assign #(out_delay) CFGFUNCTIONPOWERSTATE_OUT = delay_CFGFUNCTIONPOWERSTATE;
  assign #(out_delay) CFGFUNCTIONSTATUS_OUT = delay_CFGFUNCTIONSTATUS;
  assign #(out_delay) CFGHOTRESETOUT_OUT = delay_CFGHOTRESETOUT;
  assign #(out_delay) CFGINPUTUPDATEDONE_OUT = delay_CFGINPUTUPDATEDONE;
  assign #(out_delay) CFGINTERRUPTAOUTPUT_OUT = delay_CFGINTERRUPTAOUTPUT;
  assign #(out_delay) CFGINTERRUPTBOUTPUT_OUT = delay_CFGINTERRUPTBOUTPUT;
  assign #(out_delay) CFGINTERRUPTCOUTPUT_OUT = delay_CFGINTERRUPTCOUTPUT;
  assign #(out_delay) CFGINTERRUPTDOUTPUT_OUT = delay_CFGINTERRUPTDOUTPUT;
  assign #(out_delay) CFGINTERRUPTMSIDATA_OUT = delay_CFGINTERRUPTMSIDATA;
  assign #(out_delay) CFGINTERRUPTMSIENABLE_OUT = delay_CFGINTERRUPTMSIENABLE;
  assign #(out_delay) CFGINTERRUPTMSIFAIL_OUT = delay_CFGINTERRUPTMSIFAIL;
  assign #(out_delay) CFGINTERRUPTMSIMASKUPDATE_OUT = delay_CFGINTERRUPTMSIMASKUPDATE;
  assign #(out_delay) CFGINTERRUPTMSIMMENABLE_OUT = delay_CFGINTERRUPTMSIMMENABLE;
  assign #(out_delay) CFGINTERRUPTMSISENT_OUT = delay_CFGINTERRUPTMSISENT;
  assign #(out_delay) CFGINTERRUPTMSIVFENABLE_OUT = delay_CFGINTERRUPTMSIVFENABLE;
  assign #(out_delay) CFGINTERRUPTMSIXENABLE_OUT = delay_CFGINTERRUPTMSIXENABLE;
  assign #(out_delay) CFGINTERRUPTMSIXFAIL_OUT = delay_CFGINTERRUPTMSIXFAIL;
  assign #(out_delay) CFGINTERRUPTMSIXMASK_OUT = delay_CFGINTERRUPTMSIXMASK;
  assign #(out_delay) CFGINTERRUPTMSIXSENT_OUT = delay_CFGINTERRUPTMSIXSENT;
  assign #(out_delay) CFGINTERRUPTMSIXVFENABLE_OUT = delay_CFGINTERRUPTMSIXVFENABLE;
  assign #(out_delay) CFGINTERRUPTMSIXVFMASK_OUT = delay_CFGINTERRUPTMSIXVFMASK;
  assign #(out_delay) CFGINTERRUPTSENT_OUT = delay_CFGINTERRUPTSENT;
  assign #(out_delay) CFGLINKPOWERSTATE_OUT = delay_CFGLINKPOWERSTATE;
  assign #(out_delay) CFGLOCALERROR_OUT = delay_CFGLOCALERROR;
  assign #(out_delay) CFGLTRENABLE_OUT = delay_CFGLTRENABLE;
  assign #(out_delay) CFGLTSSMSTATE_OUT = delay_CFGLTSSMSTATE;
  assign #(out_delay) CFGMAXPAYLOAD_OUT = delay_CFGMAXPAYLOAD;
  assign #(out_delay) CFGMAXREADREQ_OUT = delay_CFGMAXREADREQ;
  assign #(out_delay) CFGMCUPDATEDONE_OUT = delay_CFGMCUPDATEDONE;
  assign #(out_delay) CFGMGMTREADDATA_OUT = delay_CFGMGMTREADDATA;
  assign #(out_delay) CFGMGMTREADWRITEDONE_OUT = delay_CFGMGMTREADWRITEDONE;
  assign #(out_delay) CFGMSGRECEIVEDDATA_OUT = delay_CFGMSGRECEIVEDDATA;
  assign #(out_delay) CFGMSGRECEIVEDTYPE_OUT = delay_CFGMSGRECEIVEDTYPE;
  assign #(out_delay) CFGMSGRECEIVED_OUT = delay_CFGMSGRECEIVED;
  assign #(out_delay) CFGMSGTRANSMITDONE_OUT = delay_CFGMSGTRANSMITDONE;
  assign #(out_delay) CFGNEGOTIATEDWIDTH_OUT = delay_CFGNEGOTIATEDWIDTH;
  assign #(out_delay) CFGOBFFENABLE_OUT = delay_CFGOBFFENABLE;
  assign #(out_delay) CFGPERFUNCSTATUSDATA_OUT = delay_CFGPERFUNCSTATUSDATA;
  assign #(out_delay) CFGPERFUNCTIONUPDATEDONE_OUT = delay_CFGPERFUNCTIONUPDATEDONE;
  assign #(out_delay) CFGPHYLINKDOWN_OUT = delay_CFGPHYLINKDOWN;
  assign #(out_delay) CFGPHYLINKSTATUS_OUT = delay_CFGPHYLINKSTATUS;
  assign #(out_delay) CFGPLSTATUSCHANGE_OUT = delay_CFGPLSTATUSCHANGE;
  assign #(out_delay) CFGPOWERSTATECHANGEINTERRUPT_OUT = delay_CFGPOWERSTATECHANGEINTERRUPT;
  assign #(out_delay) CFGRCBSTATUS_OUT = delay_CFGRCBSTATUS;
  assign #(out_delay) CFGTPHFUNCTIONNUM_OUT = delay_CFGTPHFUNCTIONNUM;
  assign #(out_delay) CFGTPHREQUESTERENABLE_OUT = delay_CFGTPHREQUESTERENABLE;
  assign #(out_delay) CFGTPHSTMODE_OUT = delay_CFGTPHSTMODE;
  assign #(out_delay) CFGTPHSTTADDRESS_OUT = delay_CFGTPHSTTADDRESS;
  assign #(out_delay) CFGTPHSTTREADENABLE_OUT = delay_CFGTPHSTTREADENABLE;
  assign #(out_delay) CFGTPHSTTWRITEBYTEVALID_OUT = delay_CFGTPHSTTWRITEBYTEVALID;
  assign #(out_delay) CFGTPHSTTWRITEDATA_OUT = delay_CFGTPHSTTWRITEDATA;
  assign #(out_delay) CFGTPHSTTWRITEENABLE_OUT = delay_CFGTPHSTTWRITEENABLE;
  assign #(out_delay) CFGVFFLRINPROCESS_OUT = delay_CFGVFFLRINPROCESS;
  assign #(out_delay) CFGVFPOWERSTATE_OUT = delay_CFGVFPOWERSTATE;
  assign #(out_delay) CFGVFSTATUS_OUT = delay_CFGVFSTATUS;
  assign #(out_delay) CFGVFTPHREQUESTERENABLE_OUT = delay_CFGVFTPHREQUESTERENABLE;
  assign #(out_delay) CFGVFTPHSTMODE_OUT = delay_CFGVFTPHSTMODE;
  assign #(out_delay) DBGDATAOUT_OUT = delay_DBGDATAOUT;
  assign #(out_delay) DRPDO_OUT = delay_DRPDO;
  assign #(out_delay) DRPRDY_OUT = delay_DRPRDY;
  assign #(out_delay) MAXISCQTDATA_OUT = delay_MAXISCQTDATA;
  assign #(out_delay) MAXISCQTKEEP_OUT = delay_MAXISCQTKEEP;
  assign #(out_delay) MAXISCQTLAST_OUT = delay_MAXISCQTLAST;
  assign #(out_delay) MAXISCQTUSER_OUT = delay_MAXISCQTUSER;
  assign #(out_delay) MAXISCQTVALID_OUT = delay_MAXISCQTVALID;
  assign #(out_delay) MAXISRCTDATA_OUT = delay_MAXISRCTDATA;
  assign #(out_delay) MAXISRCTKEEP_OUT = delay_MAXISRCTKEEP;
  assign #(out_delay) MAXISRCTLAST_OUT = delay_MAXISRCTLAST;
  assign #(out_delay) MAXISRCTUSER_OUT = delay_MAXISRCTUSER;
  assign #(out_delay) MAXISRCTVALID_OUT = delay_MAXISRCTVALID;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSAL_OUT = delay_MICOMPLETIONRAMREADADDRESSAL;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSAU_OUT = delay_MICOMPLETIONRAMREADADDRESSAU;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSBL_OUT = delay_MICOMPLETIONRAMREADADDRESSBL;
  assign #(out_delay) MICOMPLETIONRAMREADADDRESSBU_OUT = delay_MICOMPLETIONRAMREADADDRESSBU;
  assign #(out_delay) MICOMPLETIONRAMREADENABLEL_OUT = delay_MICOMPLETIONRAMREADENABLEL;
  assign #(out_delay) MICOMPLETIONRAMREADENABLEU_OUT = delay_MICOMPLETIONRAMREADENABLEU;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSAL_OUT = delay_MICOMPLETIONRAMWRITEADDRESSAL;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSAU_OUT = delay_MICOMPLETIONRAMWRITEADDRESSAU;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSBL_OUT = delay_MICOMPLETIONRAMWRITEADDRESSBL;
  assign #(out_delay) MICOMPLETIONRAMWRITEADDRESSBU_OUT = delay_MICOMPLETIONRAMWRITEADDRESSBU;
  assign #(out_delay) MICOMPLETIONRAMWRITEDATAL_OUT = delay_MICOMPLETIONRAMWRITEDATAL;
  assign #(out_delay) MICOMPLETIONRAMWRITEDATAU_OUT = delay_MICOMPLETIONRAMWRITEDATAU;
  assign #(out_delay) MICOMPLETIONRAMWRITEENABLEL_OUT = delay_MICOMPLETIONRAMWRITEENABLEL;
  assign #(out_delay) MICOMPLETIONRAMWRITEENABLEU_OUT = delay_MICOMPLETIONRAMWRITEENABLEU;
  assign #(out_delay) MIREPLAYRAMADDRESS_OUT = delay_MIREPLAYRAMADDRESS;
  assign #(out_delay) MIREPLAYRAMREADENABLE_OUT = delay_MIREPLAYRAMREADENABLE;
  assign #(out_delay) MIREPLAYRAMWRITEDATA_OUT = delay_MIREPLAYRAMWRITEDATA;
  assign #(out_delay) MIREPLAYRAMWRITEENABLE_OUT = delay_MIREPLAYRAMWRITEENABLE;
  assign #(out_delay) MIREQUESTRAMREADADDRESSA_OUT = delay_MIREQUESTRAMREADADDRESSA;
  assign #(out_delay) MIREQUESTRAMREADADDRESSB_OUT = delay_MIREQUESTRAMREADADDRESSB;
  assign #(out_delay) MIREQUESTRAMREADENABLE_OUT = delay_MIREQUESTRAMREADENABLE;
  assign #(out_delay) MIREQUESTRAMWRITEADDRESSA_OUT = delay_MIREQUESTRAMWRITEADDRESSA;
  assign #(out_delay) MIREQUESTRAMWRITEADDRESSB_OUT = delay_MIREQUESTRAMWRITEADDRESSB;
  assign #(out_delay) MIREQUESTRAMWRITEDATA_OUT = delay_MIREQUESTRAMWRITEDATA;
  assign #(out_delay) MIREQUESTRAMWRITEENABLE_OUT = delay_MIREQUESTRAMWRITEENABLE;
  assign #(out_delay) PCIECQNPREQCOUNT_OUT = delay_PCIECQNPREQCOUNT;
  assign #(out_delay) PCIERQSEQNUMVLD_OUT = delay_PCIERQSEQNUMVLD;
  assign #(out_delay) PCIERQSEQNUM_OUT = delay_PCIERQSEQNUM;
  assign #(out_delay) PCIERQTAGAV_OUT = delay_PCIERQTAGAV;
  assign #(out_delay) PCIERQTAGVLD_OUT = delay_PCIERQTAGVLD;
  assign #(out_delay) PCIERQTAG_OUT = delay_PCIERQTAG;
  assign #(out_delay) PCIETFCNPDAV_OUT = delay_PCIETFCNPDAV;
  assign #(out_delay) PCIETFCNPHAV_OUT = delay_PCIETFCNPHAV;
  assign #(out_delay) PIPERX0EQCONTROL_OUT = delay_PIPERX0EQCONTROL;
  assign #(out_delay) PIPERX0EQLPLFFS_OUT = delay_PIPERX0EQLPLFFS;
  assign #(out_delay) PIPERX0EQLPTXPRESET_OUT = delay_PIPERX0EQLPTXPRESET;
  assign #(out_delay) PIPERX0EQPRESET_OUT = delay_PIPERX0EQPRESET;
  assign #(out_delay) PIPERX0POLARITY_OUT = delay_PIPERX0POLARITY;
  assign #(out_delay) PIPERX1EQCONTROL_OUT = delay_PIPERX1EQCONTROL;
  assign #(out_delay) PIPERX1EQLPLFFS_OUT = delay_PIPERX1EQLPLFFS;
  assign #(out_delay) PIPERX1EQLPTXPRESET_OUT = delay_PIPERX1EQLPTXPRESET;
  assign #(out_delay) PIPERX1EQPRESET_OUT = delay_PIPERX1EQPRESET;
  assign #(out_delay) PIPERX1POLARITY_OUT = delay_PIPERX1POLARITY;
  assign #(out_delay) PIPERX2EQCONTROL_OUT = delay_PIPERX2EQCONTROL;
  assign #(out_delay) PIPERX2EQLPLFFS_OUT = delay_PIPERX2EQLPLFFS;
  assign #(out_delay) PIPERX2EQLPTXPRESET_OUT = delay_PIPERX2EQLPTXPRESET;
  assign #(out_delay) PIPERX2EQPRESET_OUT = delay_PIPERX2EQPRESET;
  assign #(out_delay) PIPERX2POLARITY_OUT = delay_PIPERX2POLARITY;
  assign #(out_delay) PIPERX3EQCONTROL_OUT = delay_PIPERX3EQCONTROL;
  assign #(out_delay) PIPERX3EQLPLFFS_OUT = delay_PIPERX3EQLPLFFS;
  assign #(out_delay) PIPERX3EQLPTXPRESET_OUT = delay_PIPERX3EQLPTXPRESET;
  assign #(out_delay) PIPERX3EQPRESET_OUT = delay_PIPERX3EQPRESET;
  assign #(out_delay) PIPERX3POLARITY_OUT = delay_PIPERX3POLARITY;
  assign #(out_delay) PIPERX4EQCONTROL_OUT = delay_PIPERX4EQCONTROL;
  assign #(out_delay) PIPERX4EQLPLFFS_OUT = delay_PIPERX4EQLPLFFS;
  assign #(out_delay) PIPERX4EQLPTXPRESET_OUT = delay_PIPERX4EQLPTXPRESET;
  assign #(out_delay) PIPERX4EQPRESET_OUT = delay_PIPERX4EQPRESET;
  assign #(out_delay) PIPERX4POLARITY_OUT = delay_PIPERX4POLARITY;
  assign #(out_delay) PIPERX5EQCONTROL_OUT = delay_PIPERX5EQCONTROL;
  assign #(out_delay) PIPERX5EQLPLFFS_OUT = delay_PIPERX5EQLPLFFS;
  assign #(out_delay) PIPERX5EQLPTXPRESET_OUT = delay_PIPERX5EQLPTXPRESET;
  assign #(out_delay) PIPERX5EQPRESET_OUT = delay_PIPERX5EQPRESET;
  assign #(out_delay) PIPERX5POLARITY_OUT = delay_PIPERX5POLARITY;
  assign #(out_delay) PIPERX6EQCONTROL_OUT = delay_PIPERX6EQCONTROL;
  assign #(out_delay) PIPERX6EQLPLFFS_OUT = delay_PIPERX6EQLPLFFS;
  assign #(out_delay) PIPERX6EQLPTXPRESET_OUT = delay_PIPERX6EQLPTXPRESET;
  assign #(out_delay) PIPERX6EQPRESET_OUT = delay_PIPERX6EQPRESET;
  assign #(out_delay) PIPERX6POLARITY_OUT = delay_PIPERX6POLARITY;
  assign #(out_delay) PIPERX7EQCONTROL_OUT = delay_PIPERX7EQCONTROL;
  assign #(out_delay) PIPERX7EQLPLFFS_OUT = delay_PIPERX7EQLPLFFS;
  assign #(out_delay) PIPERX7EQLPTXPRESET_OUT = delay_PIPERX7EQLPTXPRESET;
  assign #(out_delay) PIPERX7EQPRESET_OUT = delay_PIPERX7EQPRESET;
  assign #(out_delay) PIPERX7POLARITY_OUT = delay_PIPERX7POLARITY;
  assign #(out_delay) PIPETX0CHARISK_OUT = delay_PIPETX0CHARISK;
  assign #(out_delay) PIPETX0COMPLIANCE_OUT = delay_PIPETX0COMPLIANCE;
  assign #(out_delay) PIPETX0DATAVALID_OUT = delay_PIPETX0DATAVALID;
  assign #(out_delay) PIPETX0DATA_OUT = delay_PIPETX0DATA;
  assign #(out_delay) PIPETX0ELECIDLE_OUT = delay_PIPETX0ELECIDLE;
  assign #(out_delay) PIPETX0EQCONTROL_OUT = delay_PIPETX0EQCONTROL;
  assign #(out_delay) PIPETX0EQDEEMPH_OUT = delay_PIPETX0EQDEEMPH;
  assign #(out_delay) PIPETX0EQPRESET_OUT = delay_PIPETX0EQPRESET;
  assign #(out_delay) PIPETX0POWERDOWN_OUT = delay_PIPETX0POWERDOWN;
  assign #(out_delay) PIPETX0STARTBLOCK_OUT = delay_PIPETX0STARTBLOCK;
  assign #(out_delay) PIPETX0SYNCHEADER_OUT = delay_PIPETX0SYNCHEADER;
  assign #(out_delay) PIPETX1CHARISK_OUT = delay_PIPETX1CHARISK;
  assign #(out_delay) PIPETX1COMPLIANCE_OUT = delay_PIPETX1COMPLIANCE;
  assign #(out_delay) PIPETX1DATAVALID_OUT = delay_PIPETX1DATAVALID;
  assign #(out_delay) PIPETX1DATA_OUT = delay_PIPETX1DATA;
  assign #(out_delay) PIPETX1ELECIDLE_OUT = delay_PIPETX1ELECIDLE;
  assign #(out_delay) PIPETX1EQCONTROL_OUT = delay_PIPETX1EQCONTROL;
  assign #(out_delay) PIPETX1EQDEEMPH_OUT = delay_PIPETX1EQDEEMPH;
  assign #(out_delay) PIPETX1EQPRESET_OUT = delay_PIPETX1EQPRESET;
  assign #(out_delay) PIPETX1POWERDOWN_OUT = delay_PIPETX1POWERDOWN;
  assign #(out_delay) PIPETX1STARTBLOCK_OUT = delay_PIPETX1STARTBLOCK;
  assign #(out_delay) PIPETX1SYNCHEADER_OUT = delay_PIPETX1SYNCHEADER;
  assign #(out_delay) PIPETX2CHARISK_OUT = delay_PIPETX2CHARISK;
  assign #(out_delay) PIPETX2COMPLIANCE_OUT = delay_PIPETX2COMPLIANCE;
  assign #(out_delay) PIPETX2DATAVALID_OUT = delay_PIPETX2DATAVALID;
  assign #(out_delay) PIPETX2DATA_OUT = delay_PIPETX2DATA;
  assign #(out_delay) PIPETX2ELECIDLE_OUT = delay_PIPETX2ELECIDLE;
  assign #(out_delay) PIPETX2EQCONTROL_OUT = delay_PIPETX2EQCONTROL;
  assign #(out_delay) PIPETX2EQDEEMPH_OUT = delay_PIPETX2EQDEEMPH;
  assign #(out_delay) PIPETX2EQPRESET_OUT = delay_PIPETX2EQPRESET;
  assign #(out_delay) PIPETX2POWERDOWN_OUT = delay_PIPETX2POWERDOWN;
  assign #(out_delay) PIPETX2STARTBLOCK_OUT = delay_PIPETX2STARTBLOCK;
  assign #(out_delay) PIPETX2SYNCHEADER_OUT = delay_PIPETX2SYNCHEADER;
  assign #(out_delay) PIPETX3CHARISK_OUT = delay_PIPETX3CHARISK;
  assign #(out_delay) PIPETX3COMPLIANCE_OUT = delay_PIPETX3COMPLIANCE;
  assign #(out_delay) PIPETX3DATAVALID_OUT = delay_PIPETX3DATAVALID;
  assign #(out_delay) PIPETX3DATA_OUT = delay_PIPETX3DATA;
  assign #(out_delay) PIPETX3ELECIDLE_OUT = delay_PIPETX3ELECIDLE;
  assign #(out_delay) PIPETX3EQCONTROL_OUT = delay_PIPETX3EQCONTROL;
  assign #(out_delay) PIPETX3EQDEEMPH_OUT = delay_PIPETX3EQDEEMPH;
  assign #(out_delay) PIPETX3EQPRESET_OUT = delay_PIPETX3EQPRESET;
  assign #(out_delay) PIPETX3POWERDOWN_OUT = delay_PIPETX3POWERDOWN;
  assign #(out_delay) PIPETX3STARTBLOCK_OUT = delay_PIPETX3STARTBLOCK;
  assign #(out_delay) PIPETX3SYNCHEADER_OUT = delay_PIPETX3SYNCHEADER;
  assign #(out_delay) PIPETX4CHARISK_OUT = delay_PIPETX4CHARISK;
  assign #(out_delay) PIPETX4COMPLIANCE_OUT = delay_PIPETX4COMPLIANCE;
  assign #(out_delay) PIPETX4DATAVALID_OUT = delay_PIPETX4DATAVALID;
  assign #(out_delay) PIPETX4DATA_OUT = delay_PIPETX4DATA;
  assign #(out_delay) PIPETX4ELECIDLE_OUT = delay_PIPETX4ELECIDLE;
  assign #(out_delay) PIPETX4EQCONTROL_OUT = delay_PIPETX4EQCONTROL;
  assign #(out_delay) PIPETX4EQDEEMPH_OUT = delay_PIPETX4EQDEEMPH;
  assign #(out_delay) PIPETX4EQPRESET_OUT = delay_PIPETX4EQPRESET;
  assign #(out_delay) PIPETX4POWERDOWN_OUT = delay_PIPETX4POWERDOWN;
  assign #(out_delay) PIPETX4STARTBLOCK_OUT = delay_PIPETX4STARTBLOCK;
  assign #(out_delay) PIPETX4SYNCHEADER_OUT = delay_PIPETX4SYNCHEADER;
  assign #(out_delay) PIPETX5CHARISK_OUT = delay_PIPETX5CHARISK;
  assign #(out_delay) PIPETX5COMPLIANCE_OUT = delay_PIPETX5COMPLIANCE;
  assign #(out_delay) PIPETX5DATAVALID_OUT = delay_PIPETX5DATAVALID;
  assign #(out_delay) PIPETX5DATA_OUT = delay_PIPETX5DATA;
  assign #(out_delay) PIPETX5ELECIDLE_OUT = delay_PIPETX5ELECIDLE;
  assign #(out_delay) PIPETX5EQCONTROL_OUT = delay_PIPETX5EQCONTROL;
  assign #(out_delay) PIPETX5EQDEEMPH_OUT = delay_PIPETX5EQDEEMPH;
  assign #(out_delay) PIPETX5EQPRESET_OUT = delay_PIPETX5EQPRESET;
  assign #(out_delay) PIPETX5POWERDOWN_OUT = delay_PIPETX5POWERDOWN;
  assign #(out_delay) PIPETX5STARTBLOCK_OUT = delay_PIPETX5STARTBLOCK;
  assign #(out_delay) PIPETX5SYNCHEADER_OUT = delay_PIPETX5SYNCHEADER;
  assign #(out_delay) PIPETX6CHARISK_OUT = delay_PIPETX6CHARISK;
  assign #(out_delay) PIPETX6COMPLIANCE_OUT = delay_PIPETX6COMPLIANCE;
  assign #(out_delay) PIPETX6DATAVALID_OUT = delay_PIPETX6DATAVALID;
  assign #(out_delay) PIPETX6DATA_OUT = delay_PIPETX6DATA;
  assign #(out_delay) PIPETX6ELECIDLE_OUT = delay_PIPETX6ELECIDLE;
  assign #(out_delay) PIPETX6EQCONTROL_OUT = delay_PIPETX6EQCONTROL;
  assign #(out_delay) PIPETX6EQDEEMPH_OUT = delay_PIPETX6EQDEEMPH;
  assign #(out_delay) PIPETX6EQPRESET_OUT = delay_PIPETX6EQPRESET;
  assign #(out_delay) PIPETX6POWERDOWN_OUT = delay_PIPETX6POWERDOWN;
  assign #(out_delay) PIPETX6STARTBLOCK_OUT = delay_PIPETX6STARTBLOCK;
  assign #(out_delay) PIPETX6SYNCHEADER_OUT = delay_PIPETX6SYNCHEADER;
  assign #(out_delay) PIPETX7CHARISK_OUT = delay_PIPETX7CHARISK;
  assign #(out_delay) PIPETX7COMPLIANCE_OUT = delay_PIPETX7COMPLIANCE;
  assign #(out_delay) PIPETX7DATAVALID_OUT = delay_PIPETX7DATAVALID;
  assign #(out_delay) PIPETX7DATA_OUT = delay_PIPETX7DATA;
  assign #(out_delay) PIPETX7ELECIDLE_OUT = delay_PIPETX7ELECIDLE;
  assign #(out_delay) PIPETX7EQCONTROL_OUT = delay_PIPETX7EQCONTROL;
  assign #(out_delay) PIPETX7EQDEEMPH_OUT = delay_PIPETX7EQDEEMPH;
  assign #(out_delay) PIPETX7EQPRESET_OUT = delay_PIPETX7EQPRESET;
  assign #(out_delay) PIPETX7POWERDOWN_OUT = delay_PIPETX7POWERDOWN;
  assign #(out_delay) PIPETX7STARTBLOCK_OUT = delay_PIPETX7STARTBLOCK;
  assign #(out_delay) PIPETX7SYNCHEADER_OUT = delay_PIPETX7SYNCHEADER;
  assign #(out_delay) PIPETXDEEMPH_OUT = delay_PIPETXDEEMPH;
  assign #(out_delay) PIPETXMARGIN_OUT = delay_PIPETXMARGIN;
  assign #(out_delay) PIPETXRATE_OUT = delay_PIPETXRATE;
  assign #(out_delay) PIPETXRCVRDET_OUT = delay_PIPETXRCVRDET;
  assign #(out_delay) PIPETXRESET_OUT = delay_PIPETXRESET;
  assign #(out_delay) PIPETXSWING_OUT = delay_PIPETXSWING;
  assign #(out_delay) PLEQINPROGRESS_OUT = delay_PLEQINPROGRESS;
  assign #(out_delay) PLEQPHASE_OUT = delay_PLEQPHASE;
  assign #(out_delay) PLGEN3PCSRXSLIDE_OUT = delay_PLGEN3PCSRXSLIDE;
  assign #(out_delay) SAXISCCTREADY_OUT = delay_SAXISCCTREADY;
  assign #(out_delay) SAXISRQTREADY_OUT = delay_SAXISRQTREADY;

  assign #(INCLK_DELAY) CORECLKMICOMPLETIONRAML_INDELAY = CORECLKMICOMPLETIONRAML_IN;
  assign #(INCLK_DELAY) CORECLKMICOMPLETIONRAMU_INDELAY = CORECLKMICOMPLETIONRAMU_IN;
  assign #(INCLK_DELAY) CORECLKMIREPLAYRAM_INDELAY = CORECLKMIREPLAYRAM_IN;
  assign #(INCLK_DELAY) CORECLKMIREQUESTRAM_INDELAY = CORECLKMIREQUESTRAM_IN;
  assign #(INCLK_DELAY) CORECLK_INDELAY = CORECLK_IN;
  assign #(INCLK_DELAY) DRPCLK_INDELAY = DRPCLK_IN;
  assign #(INCLK_DELAY) PIPECLK_INDELAY = PIPECLK_IN;
  assign #(INCLK_DELAY) RECCLK_INDELAY = RECCLK_IN;
  assign #(INCLK_DELAY) USERCLK_INDELAY = USERCLK_IN;

  assign #(in_delay) CFGCONFIGSPACEENABLE_INDELAY = CFGCONFIGSPACEENABLE_IN;
  assign #(in_delay) CFGDEVID_INDELAY = CFGDEVID_IN;
  assign #(in_delay) CFGDSBUSNUMBER_INDELAY = CFGDSBUSNUMBER_IN;
  assign #(in_delay) CFGDSDEVICENUMBER_INDELAY = CFGDSDEVICENUMBER_IN;
  assign #(in_delay) CFGDSFUNCTIONNUMBER_INDELAY = CFGDSFUNCTIONNUMBER_IN;
  assign #(in_delay) CFGDSN_INDELAY = CFGDSN_IN;
  assign #(in_delay) CFGDSPORTNUMBER_INDELAY = CFGDSPORTNUMBER_IN;
  assign #(in_delay) CFGERRCORIN_INDELAY = CFGERRCORIN_IN;
  assign #(in_delay) CFGERRUNCORIN_INDELAY = CFGERRUNCORIN_IN;
  assign #(in_delay) CFGEXTREADDATAVALID_INDELAY = CFGEXTREADDATAVALID_IN;
  assign #(in_delay) CFGEXTREADDATA_INDELAY = CFGEXTREADDATA_IN;
  assign #(in_delay) CFGFCSEL_INDELAY = CFGFCSEL_IN;
  assign #(in_delay) CFGFLRDONE_INDELAY = CFGFLRDONE_IN;
  assign #(in_delay) CFGHOTRESETIN_INDELAY = CFGHOTRESETIN_IN;
  assign #(in_delay) CFGINPUTUPDATEREQUEST_INDELAY = CFGINPUTUPDATEREQUEST_IN;
  assign #(in_delay) CFGINTERRUPTINT_INDELAY = CFGINTERRUPTINT_IN;
  assign #(in_delay) CFGINTERRUPTMSIATTR_INDELAY = CFGINTERRUPTMSIATTR_IN;
  assign #(in_delay) CFGINTERRUPTMSIFUNCTIONNUMBER_INDELAY = CFGINTERRUPTMSIFUNCTIONNUMBER_IN;
  assign #(in_delay) CFGINTERRUPTMSIINT_INDELAY = CFGINTERRUPTMSIINT_IN;
  assign #(in_delay) CFGINTERRUPTMSIPENDINGSTATUS_INDELAY = CFGINTERRUPTMSIPENDINGSTATUS_IN;
  assign #(in_delay) CFGINTERRUPTMSISELECT_INDELAY = CFGINTERRUPTMSISELECT_IN;
  assign #(in_delay) CFGINTERRUPTMSITPHPRESENT_INDELAY = CFGINTERRUPTMSITPHPRESENT_IN;
  assign #(in_delay) CFGINTERRUPTMSITPHSTTAG_INDELAY = CFGINTERRUPTMSITPHSTTAG_IN;
  assign #(in_delay) CFGINTERRUPTMSITPHTYPE_INDELAY = CFGINTERRUPTMSITPHTYPE_IN;
  assign #(in_delay) CFGINTERRUPTMSIXADDRESS_INDELAY = CFGINTERRUPTMSIXADDRESS_IN;
  assign #(in_delay) CFGINTERRUPTMSIXDATA_INDELAY = CFGINTERRUPTMSIXDATA_IN;
  assign #(in_delay) CFGINTERRUPTMSIXINT_INDELAY = CFGINTERRUPTMSIXINT_IN;
  assign #(in_delay) CFGINTERRUPTPENDING_INDELAY = CFGINTERRUPTPENDING_IN;
  assign #(in_delay) CFGLINKTRAININGENABLE_INDELAY = CFGLINKTRAININGENABLE_IN;
  assign #(in_delay) CFGMCUPDATEREQUEST_INDELAY = CFGMCUPDATEREQUEST_IN;
  assign #(in_delay) CFGMGMTADDR_INDELAY = CFGMGMTADDR_IN;
  assign #(in_delay) CFGMGMTBYTEENABLE_INDELAY = CFGMGMTBYTEENABLE_IN;
  assign #(in_delay) CFGMGMTREAD_INDELAY = CFGMGMTREAD_IN;
  assign #(in_delay) CFGMGMTTYPE1CFGREGACCESS_INDELAY = CFGMGMTTYPE1CFGREGACCESS_IN;
  assign #(in_delay) CFGMGMTWRITEDATA_INDELAY = CFGMGMTWRITEDATA_IN;
  assign #(in_delay) CFGMGMTWRITE_INDELAY = CFGMGMTWRITE_IN;
  assign #(in_delay) CFGMSGTRANSMITDATA_INDELAY = CFGMSGTRANSMITDATA_IN;
  assign #(in_delay) CFGMSGTRANSMITTYPE_INDELAY = CFGMSGTRANSMITTYPE_IN;
  assign #(in_delay) CFGMSGTRANSMIT_INDELAY = CFGMSGTRANSMIT_IN;
  assign #(in_delay) CFGPERFUNCSTATUSCONTROL_INDELAY = CFGPERFUNCSTATUSCONTROL_IN;
  assign #(in_delay) CFGPERFUNCTIONNUMBER_INDELAY = CFGPERFUNCTIONNUMBER_IN;
  assign #(in_delay) CFGPERFUNCTIONOUTPUTREQUEST_INDELAY = CFGPERFUNCTIONOUTPUTREQUEST_IN;
  assign #(in_delay) CFGPOWERSTATECHANGEACK_INDELAY = CFGPOWERSTATECHANGEACK_IN;
  assign #(in_delay) CFGREQPMTRANSITIONL23READY_INDELAY = CFGREQPMTRANSITIONL23READY_IN;
  assign #(in_delay) CFGREVID_INDELAY = CFGREVID_IN;
  assign #(in_delay) CFGSUBSYSID_INDELAY = CFGSUBSYSID_IN;
  assign #(in_delay) CFGSUBSYSVENDID_INDELAY = CFGSUBSYSVENDID_IN;
  assign #(in_delay) CFGTPHSTTREADDATAVALID_INDELAY = CFGTPHSTTREADDATAVALID_IN;
  assign #(in_delay) CFGTPHSTTREADDATA_INDELAY = CFGTPHSTTREADDATA_IN;
  assign #(in_delay) CFGVENDID_INDELAY = CFGVENDID_IN;
  assign #(in_delay) CFGVFFLRDONE_INDELAY = CFGVFFLRDONE_IN;
  assign #(in_delay) DRPADDR_INDELAY = DRPADDR_IN;
  assign #(in_delay) DRPDI_INDELAY = DRPDI_IN;
  assign #(in_delay) DRPEN_INDELAY = DRPEN_IN;
  assign #(in_delay) DRPWE_INDELAY = DRPWE_IN;
  assign #(in_delay) MAXISCQTREADY_INDELAY = MAXISCQTREADY_IN;
  assign #(in_delay) MAXISRCTREADY_INDELAY = MAXISRCTREADY_IN;
  assign #(in_delay) MGMTRESETN_INDELAY = MGMTRESETN_IN;
  assign #(in_delay) MGMTSTICKYRESETN_INDELAY = MGMTSTICKYRESETN_IN;
  assign #(in_delay) MICOMPLETIONRAMREADDATA_INDELAY = MICOMPLETIONRAMREADDATA_IN;
  assign #(in_delay) MIREPLAYRAMREADDATA_INDELAY = MIREPLAYRAMREADDATA_IN;
  assign #(in_delay) MIREQUESTRAMREADDATA_INDELAY = MIREQUESTRAMREADDATA_IN;
  assign #(in_delay) PCIECQNPREQ_INDELAY = PCIECQNPREQ_IN;
  assign #(in_delay) PIPEEQFS_INDELAY = PIPEEQFS_IN;
  assign #(in_delay) PIPEEQLF_INDELAY = PIPEEQLF_IN;
  assign #(in_delay) PIPERESETN_INDELAY = PIPERESETN_IN;
  assign #(in_delay) PIPERX0CHARISK_INDELAY = PIPERX0CHARISK_IN;
  assign #(in_delay) PIPERX0DATAVALID_INDELAY = PIPERX0DATAVALID_IN;
  assign #(in_delay) PIPERX0DATA_INDELAY = PIPERX0DATA_IN;
  assign #(in_delay) PIPERX0ELECIDLE_INDELAY = PIPERX0ELECIDLE_IN;
  assign #(in_delay) PIPERX0EQDONE_INDELAY = PIPERX0EQDONE_IN;
  assign #(in_delay) PIPERX0EQLPADAPTDONE_INDELAY = PIPERX0EQLPADAPTDONE_IN;
  assign #(in_delay) PIPERX0EQLPLFFSSEL_INDELAY = PIPERX0EQLPLFFSSEL_IN;
  assign #(in_delay) PIPERX0EQLPNEWTXCOEFFORPRESET_INDELAY = PIPERX0EQLPNEWTXCOEFFORPRESET_IN;
  assign #(in_delay) PIPERX0PHYSTATUS_INDELAY = PIPERX0PHYSTATUS_IN;
  assign #(in_delay) PIPERX0STARTBLOCK_INDELAY = PIPERX0STARTBLOCK_IN;
  assign #(in_delay) PIPERX0STATUS_INDELAY = PIPERX0STATUS_IN;
  assign #(in_delay) PIPERX0SYNCHEADER_INDELAY = PIPERX0SYNCHEADER_IN;
  assign #(in_delay) PIPERX0VALID_INDELAY = PIPERX0VALID_IN;
  assign #(in_delay) PIPERX1CHARISK_INDELAY = PIPERX1CHARISK_IN;
  assign #(in_delay) PIPERX1DATAVALID_INDELAY = PIPERX1DATAVALID_IN;
  assign #(in_delay) PIPERX1DATA_INDELAY = PIPERX1DATA_IN;
  assign #(in_delay) PIPERX1ELECIDLE_INDELAY = PIPERX1ELECIDLE_IN;
  assign #(in_delay) PIPERX1EQDONE_INDELAY = PIPERX1EQDONE_IN;
  assign #(in_delay) PIPERX1EQLPADAPTDONE_INDELAY = PIPERX1EQLPADAPTDONE_IN;
  assign #(in_delay) PIPERX1EQLPLFFSSEL_INDELAY = PIPERX1EQLPLFFSSEL_IN;
  assign #(in_delay) PIPERX1EQLPNEWTXCOEFFORPRESET_INDELAY = PIPERX1EQLPNEWTXCOEFFORPRESET_IN;
  assign #(in_delay) PIPERX1PHYSTATUS_INDELAY = PIPERX1PHYSTATUS_IN;
  assign #(in_delay) PIPERX1STARTBLOCK_INDELAY = PIPERX1STARTBLOCK_IN;
  assign #(in_delay) PIPERX1STATUS_INDELAY = PIPERX1STATUS_IN;
  assign #(in_delay) PIPERX1SYNCHEADER_INDELAY = PIPERX1SYNCHEADER_IN;
  assign #(in_delay) PIPERX1VALID_INDELAY = PIPERX1VALID_IN;
  assign #(in_delay) PIPERX2CHARISK_INDELAY = PIPERX2CHARISK_IN;
  assign #(in_delay) PIPERX2DATAVALID_INDELAY = PIPERX2DATAVALID_IN;
  assign #(in_delay) PIPERX2DATA_INDELAY = PIPERX2DATA_IN;
  assign #(in_delay) PIPERX2ELECIDLE_INDELAY = PIPERX2ELECIDLE_IN;
  assign #(in_delay) PIPERX2EQDONE_INDELAY = PIPERX2EQDONE_IN;
  assign #(in_delay) PIPERX2EQLPADAPTDONE_INDELAY = PIPERX2EQLPADAPTDONE_IN;
  assign #(in_delay) PIPERX2EQLPLFFSSEL_INDELAY = PIPERX2EQLPLFFSSEL_IN;
  assign #(in_delay) PIPERX2EQLPNEWTXCOEFFORPRESET_INDELAY = PIPERX2EQLPNEWTXCOEFFORPRESET_IN;
  assign #(in_delay) PIPERX2PHYSTATUS_INDELAY = PIPERX2PHYSTATUS_IN;
  assign #(in_delay) PIPERX2STARTBLOCK_INDELAY = PIPERX2STARTBLOCK_IN;
  assign #(in_delay) PIPERX2STATUS_INDELAY = PIPERX2STATUS_IN;
  assign #(in_delay) PIPERX2SYNCHEADER_INDELAY = PIPERX2SYNCHEADER_IN;
  assign #(in_delay) PIPERX2VALID_INDELAY = PIPERX2VALID_IN;
  assign #(in_delay) PIPERX3CHARISK_INDELAY = PIPERX3CHARISK_IN;
  assign #(in_delay) PIPERX3DATAVALID_INDELAY = PIPERX3DATAVALID_IN;
  assign #(in_delay) PIPERX3DATA_INDELAY = PIPERX3DATA_IN;
  assign #(in_delay) PIPERX3ELECIDLE_INDELAY = PIPERX3ELECIDLE_IN;
  assign #(in_delay) PIPERX3EQDONE_INDELAY = PIPERX3EQDONE_IN;
  assign #(in_delay) PIPERX3EQLPADAPTDONE_INDELAY = PIPERX3EQLPADAPTDONE_IN;
  assign #(in_delay) PIPERX3EQLPLFFSSEL_INDELAY = PIPERX3EQLPLFFSSEL_IN;
  assign #(in_delay) PIPERX3EQLPNEWTXCOEFFORPRESET_INDELAY = PIPERX3EQLPNEWTXCOEFFORPRESET_IN;
  assign #(in_delay) PIPERX3PHYSTATUS_INDELAY = PIPERX3PHYSTATUS_IN;
  assign #(in_delay) PIPERX3STARTBLOCK_INDELAY = PIPERX3STARTBLOCK_IN;
  assign #(in_delay) PIPERX3STATUS_INDELAY = PIPERX3STATUS_IN;
  assign #(in_delay) PIPERX3SYNCHEADER_INDELAY = PIPERX3SYNCHEADER_IN;
  assign #(in_delay) PIPERX3VALID_INDELAY = PIPERX3VALID_IN;
  assign #(in_delay) PIPERX4CHARISK_INDELAY = PIPERX4CHARISK_IN;
  assign #(in_delay) PIPERX4DATAVALID_INDELAY = PIPERX4DATAVALID_IN;
  assign #(in_delay) PIPERX4DATA_INDELAY = PIPERX4DATA_IN;
  assign #(in_delay) PIPERX4ELECIDLE_INDELAY = PIPERX4ELECIDLE_IN;
  assign #(in_delay) PIPERX4EQDONE_INDELAY = PIPERX4EQDONE_IN;
  assign #(in_delay) PIPERX4EQLPADAPTDONE_INDELAY = PIPERX4EQLPADAPTDONE_IN;
  assign #(in_delay) PIPERX4EQLPLFFSSEL_INDELAY = PIPERX4EQLPLFFSSEL_IN;
  assign #(in_delay) PIPERX4EQLPNEWTXCOEFFORPRESET_INDELAY = PIPERX4EQLPNEWTXCOEFFORPRESET_IN;
  assign #(in_delay) PIPERX4PHYSTATUS_INDELAY = PIPERX4PHYSTATUS_IN;
  assign #(in_delay) PIPERX4STARTBLOCK_INDELAY = PIPERX4STARTBLOCK_IN;
  assign #(in_delay) PIPERX4STATUS_INDELAY = PIPERX4STATUS_IN;
  assign #(in_delay) PIPERX4SYNCHEADER_INDELAY = PIPERX4SYNCHEADER_IN;
  assign #(in_delay) PIPERX4VALID_INDELAY = PIPERX4VALID_IN;
  assign #(in_delay) PIPERX5CHARISK_INDELAY = PIPERX5CHARISK_IN;
  assign #(in_delay) PIPERX5DATAVALID_INDELAY = PIPERX5DATAVALID_IN;
  assign #(in_delay) PIPERX5DATA_INDELAY = PIPERX5DATA_IN;
  assign #(in_delay) PIPERX5ELECIDLE_INDELAY = PIPERX5ELECIDLE_IN;
  assign #(in_delay) PIPERX5EQDONE_INDELAY = PIPERX5EQDONE_IN;
  assign #(in_delay) PIPERX5EQLPADAPTDONE_INDELAY = PIPERX5EQLPADAPTDONE_IN;
  assign #(in_delay) PIPERX5EQLPLFFSSEL_INDELAY = PIPERX5EQLPLFFSSEL_IN;
  assign #(in_delay) PIPERX5EQLPNEWTXCOEFFORPRESET_INDELAY = PIPERX5EQLPNEWTXCOEFFORPRESET_IN;
  assign #(in_delay) PIPERX5PHYSTATUS_INDELAY = PIPERX5PHYSTATUS_IN;
  assign #(in_delay) PIPERX5STARTBLOCK_INDELAY = PIPERX5STARTBLOCK_IN;
  assign #(in_delay) PIPERX5STATUS_INDELAY = PIPERX5STATUS_IN;
  assign #(in_delay) PIPERX5SYNCHEADER_INDELAY = PIPERX5SYNCHEADER_IN;
  assign #(in_delay) PIPERX5VALID_INDELAY = PIPERX5VALID_IN;
  assign #(in_delay) PIPERX6CHARISK_INDELAY = PIPERX6CHARISK_IN;
  assign #(in_delay) PIPERX6DATAVALID_INDELAY = PIPERX6DATAVALID_IN;
  assign #(in_delay) PIPERX6DATA_INDELAY = PIPERX6DATA_IN;
  assign #(in_delay) PIPERX6ELECIDLE_INDELAY = PIPERX6ELECIDLE_IN;
  assign #(in_delay) PIPERX6EQDONE_INDELAY = PIPERX6EQDONE_IN;
  assign #(in_delay) PIPERX6EQLPADAPTDONE_INDELAY = PIPERX6EQLPADAPTDONE_IN;
  assign #(in_delay) PIPERX6EQLPLFFSSEL_INDELAY = PIPERX6EQLPLFFSSEL_IN;
  assign #(in_delay) PIPERX6EQLPNEWTXCOEFFORPRESET_INDELAY = PIPERX6EQLPNEWTXCOEFFORPRESET_IN;
  assign #(in_delay) PIPERX6PHYSTATUS_INDELAY = PIPERX6PHYSTATUS_IN;
  assign #(in_delay) PIPERX6STARTBLOCK_INDELAY = PIPERX6STARTBLOCK_IN;
  assign #(in_delay) PIPERX6STATUS_INDELAY = PIPERX6STATUS_IN;
  assign #(in_delay) PIPERX6SYNCHEADER_INDELAY = PIPERX6SYNCHEADER_IN;
  assign #(in_delay) PIPERX6VALID_INDELAY = PIPERX6VALID_IN;
  assign #(in_delay) PIPERX7CHARISK_INDELAY = PIPERX7CHARISK_IN;
  assign #(in_delay) PIPERX7DATAVALID_INDELAY = PIPERX7DATAVALID_IN;
  assign #(in_delay) PIPERX7DATA_INDELAY = PIPERX7DATA_IN;
  assign #(in_delay) PIPERX7ELECIDLE_INDELAY = PIPERX7ELECIDLE_IN;
  assign #(in_delay) PIPERX7EQDONE_INDELAY = PIPERX7EQDONE_IN;
  assign #(in_delay) PIPERX7EQLPADAPTDONE_INDELAY = PIPERX7EQLPADAPTDONE_IN;
  assign #(in_delay) PIPERX7EQLPLFFSSEL_INDELAY = PIPERX7EQLPLFFSSEL_IN;
  assign #(in_delay) PIPERX7EQLPNEWTXCOEFFORPRESET_INDELAY = PIPERX7EQLPNEWTXCOEFFORPRESET_IN;
  assign #(in_delay) PIPERX7PHYSTATUS_INDELAY = PIPERX7PHYSTATUS_IN;
  assign #(in_delay) PIPERX7STARTBLOCK_INDELAY = PIPERX7STARTBLOCK_IN;
  assign #(in_delay) PIPERX7STATUS_INDELAY = PIPERX7STATUS_IN;
  assign #(in_delay) PIPERX7SYNCHEADER_INDELAY = PIPERX7SYNCHEADER_IN;
  assign #(in_delay) PIPERX7VALID_INDELAY = PIPERX7VALID_IN;
  assign #(in_delay) PIPETX0EQCOEFF_INDELAY = PIPETX0EQCOEFF_IN;
  assign #(in_delay) PIPETX0EQDONE_INDELAY = PIPETX0EQDONE_IN;
  assign #(in_delay) PIPETX1EQCOEFF_INDELAY = PIPETX1EQCOEFF_IN;
  assign #(in_delay) PIPETX1EQDONE_INDELAY = PIPETX1EQDONE_IN;
  assign #(in_delay) PIPETX2EQCOEFF_INDELAY = PIPETX2EQCOEFF_IN;
  assign #(in_delay) PIPETX2EQDONE_INDELAY = PIPETX2EQDONE_IN;
  assign #(in_delay) PIPETX3EQCOEFF_INDELAY = PIPETX3EQCOEFF_IN;
  assign #(in_delay) PIPETX3EQDONE_INDELAY = PIPETX3EQDONE_IN;
  assign #(in_delay) PIPETX4EQCOEFF_INDELAY = PIPETX4EQCOEFF_IN;
  assign #(in_delay) PIPETX4EQDONE_INDELAY = PIPETX4EQDONE_IN;
  assign #(in_delay) PIPETX5EQCOEFF_INDELAY = PIPETX5EQCOEFF_IN;
  assign #(in_delay) PIPETX5EQDONE_INDELAY = PIPETX5EQDONE_IN;
  assign #(in_delay) PIPETX6EQCOEFF_INDELAY = PIPETX6EQCOEFF_IN;
  assign #(in_delay) PIPETX6EQDONE_INDELAY = PIPETX6EQDONE_IN;
  assign #(in_delay) PIPETX7EQCOEFF_INDELAY = PIPETX7EQCOEFF_IN;
  assign #(in_delay) PIPETX7EQDONE_INDELAY = PIPETX7EQDONE_IN;
  assign #(in_delay) PLDISABLESCRAMBLER_INDELAY = PLDISABLESCRAMBLER_IN;
  assign #(in_delay) PLEQRESETEIEOSCOUNT_INDELAY = PLEQRESETEIEOSCOUNT_IN;
  assign #(in_delay) PLGEN3PCSDISABLE_INDELAY = PLGEN3PCSDISABLE_IN;
  assign #(in_delay) PLGEN3PCSRXSYNCDONE_INDELAY = PLGEN3PCSRXSYNCDONE_IN;
  assign #(in_delay) RESETN_INDELAY = RESETN_IN;
  assign #(in_delay) SAXISCCTDATA_INDELAY = SAXISCCTDATA_IN;
  assign #(in_delay) SAXISCCTKEEP_INDELAY = SAXISCCTKEEP_IN;
  assign #(in_delay) SAXISCCTLAST_INDELAY = SAXISCCTLAST_IN;
  assign #(in_delay) SAXISCCTUSER_INDELAY = SAXISCCTUSER_IN;
  assign #(in_delay) SAXISCCTVALID_INDELAY = SAXISCCTVALID_IN;
  assign #(in_delay) SAXISRQTDATA_INDELAY = SAXISRQTDATA_IN;
  assign #(in_delay) SAXISRQTKEEP_INDELAY = SAXISRQTKEEP_IN;
  assign #(in_delay) SAXISRQTLAST_INDELAY = SAXISRQTLAST_IN;
  assign #(in_delay) SAXISRQTUSER_INDELAY = SAXISRQTUSER_IN;
  assign #(in_delay) SAXISRQTVALID_INDELAY = SAXISRQTVALID_IN;
  assign delay_CORECLKMICOMPLETIONRAML = CORECLKMICOMPLETIONRAML_INDELAY;
  assign delay_CORECLKMICOMPLETIONRAMU = CORECLKMICOMPLETIONRAMU_INDELAY;
  assign delay_CORECLKMIREPLAYRAM = CORECLKMIREPLAYRAM_INDELAY;
  assign delay_CORECLKMIREQUESTRAM = CORECLKMIREQUESTRAM_INDELAY;
  assign delay_MGMTRESETN = MGMTRESETN_INDELAY;
  assign delay_MGMTSTICKYRESETN = MGMTSTICKYRESETN_INDELAY;
  assign delay_PIPERESETN = PIPERESETN_INDELAY;
  assign delay_RESETN = RESETN_INDELAY;

  B_PCIE_3_0 #(
    .ARI_CAP_ENABLE (ARI_CAP_ENABLE),
    .AXISTEN_IF_CC_ALIGNMENT_MODE (AXISTEN_IF_CC_ALIGNMENT_MODE),
    .AXISTEN_IF_CC_PARITY_CHK (AXISTEN_IF_CC_PARITY_CHK),
    .AXISTEN_IF_CQ_ALIGNMENT_MODE (AXISTEN_IF_CQ_ALIGNMENT_MODE),
    .AXISTEN_IF_ENABLE_CLIENT_TAG (AXISTEN_IF_ENABLE_CLIENT_TAG),
    .AXISTEN_IF_ENABLE_MSG_ROUTE (AXISTEN_IF_ENABLE_MSG_ROUTE),
    .AXISTEN_IF_ENABLE_RX_MSG_INTFC (AXISTEN_IF_ENABLE_RX_MSG_INTFC),
    .AXISTEN_IF_RC_ALIGNMENT_MODE (AXISTEN_IF_RC_ALIGNMENT_MODE),
    .AXISTEN_IF_RC_STRADDLE (AXISTEN_IF_RC_STRADDLE),
    .AXISTEN_IF_RQ_ALIGNMENT_MODE (AXISTEN_IF_RQ_ALIGNMENT_MODE),
    .AXISTEN_IF_RQ_PARITY_CHK (AXISTEN_IF_RQ_PARITY_CHK),
    .AXISTEN_IF_WIDTH (AXISTEN_IF_WIDTH),
    .CRM_CORE_CLK_FREQ_500 (CRM_CORE_CLK_FREQ_500),
    .CRM_USER_CLK_FREQ (CRM_USER_CLK_FREQ),
    .DNSTREAM_LINK_NUM (DNSTREAM_LINK_NUM),
    .GEN3_PCS_AUTO_REALIGN (GEN3_PCS_AUTO_REALIGN),
    .GEN3_PCS_RX_ELECIDLE_INTERNAL (GEN3_PCS_RX_ELECIDLE_INTERNAL),
    .LL_ACK_TIMEOUT (LL_ACK_TIMEOUT),
    .LL_ACK_TIMEOUT_EN (LL_ACK_TIMEOUT_EN),
    .LL_ACK_TIMEOUT_FUNC (LL_ACK_TIMEOUT_FUNC),
    .LL_CPL_FC_UPDATE_TIMER (LL_CPL_FC_UPDATE_TIMER),
    .LL_CPL_FC_UPDATE_TIMER_OVERRIDE (LL_CPL_FC_UPDATE_TIMER_OVERRIDE),
    .LL_FC_UPDATE_TIMER (LL_FC_UPDATE_TIMER),
    .LL_FC_UPDATE_TIMER_OVERRIDE (LL_FC_UPDATE_TIMER_OVERRIDE),
    .LL_NP_FC_UPDATE_TIMER (LL_NP_FC_UPDATE_TIMER),
    .LL_NP_FC_UPDATE_TIMER_OVERRIDE (LL_NP_FC_UPDATE_TIMER_OVERRIDE),
    .LL_P_FC_UPDATE_TIMER (LL_P_FC_UPDATE_TIMER),
    .LL_P_FC_UPDATE_TIMER_OVERRIDE (LL_P_FC_UPDATE_TIMER_OVERRIDE),
    .LL_REPLAY_TIMEOUT (LL_REPLAY_TIMEOUT),
    .LL_REPLAY_TIMEOUT_EN (LL_REPLAY_TIMEOUT_EN),
    .LL_REPLAY_TIMEOUT_FUNC (LL_REPLAY_TIMEOUT_FUNC),
    .LTR_TX_MESSAGE_MINIMUM_INTERVAL (LTR_TX_MESSAGE_MINIMUM_INTERVAL),
    .LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE (LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE),
    .LTR_TX_MESSAGE_ON_LTR_ENABLE (LTR_TX_MESSAGE_ON_LTR_ENABLE),
    .PF0_AER_CAP_ECRC_CHECK_CAPABLE (PF0_AER_CAP_ECRC_CHECK_CAPABLE),
    .PF0_AER_CAP_ECRC_GEN_CAPABLE (PF0_AER_CAP_ECRC_GEN_CAPABLE),
    .PF0_AER_CAP_NEXTPTR (PF0_AER_CAP_NEXTPTR),
    .PF0_ARI_CAP_NEXTPTR (PF0_ARI_CAP_NEXTPTR),
    .PF0_ARI_CAP_NEXT_FUNC (PF0_ARI_CAP_NEXT_FUNC),
    .PF0_ARI_CAP_VER (PF0_ARI_CAP_VER),
    .PF0_BAR0_APERTURE_SIZE (PF0_BAR0_APERTURE_SIZE),
    .PF0_BAR0_CONTROL (PF0_BAR0_CONTROL),
    .PF0_BAR1_APERTURE_SIZE (PF0_BAR1_APERTURE_SIZE),
    .PF0_BAR1_CONTROL (PF0_BAR1_CONTROL),
    .PF0_BAR2_APERTURE_SIZE (PF0_BAR2_APERTURE_SIZE),
    .PF0_BAR2_CONTROL (PF0_BAR2_CONTROL),
    .PF0_BAR3_APERTURE_SIZE (PF0_BAR3_APERTURE_SIZE),
    .PF0_BAR3_CONTROL (PF0_BAR3_CONTROL),
    .PF0_BAR4_APERTURE_SIZE (PF0_BAR4_APERTURE_SIZE),
    .PF0_BAR4_CONTROL (PF0_BAR4_CONTROL),
    .PF0_BAR5_APERTURE_SIZE (PF0_BAR5_APERTURE_SIZE),
    .PF0_BAR5_CONTROL (PF0_BAR5_CONTROL),
    .PF0_BIST_REGISTER (PF0_BIST_REGISTER),
    .PF0_CAPABILITY_POINTER (PF0_CAPABILITY_POINTER),
    .PF0_CLASS_CODE (PF0_CLASS_CODE),
    .PF0_DEVICE_ID (PF0_DEVICE_ID),
    .PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT (PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT),
    .PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT (PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT),
    .PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT (PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT),
    .PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE (PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE),
    .PF0_DEV_CAP2_LTR_SUPPORT (PF0_DEV_CAP2_LTR_SUPPORT),
    .PF0_DEV_CAP2_OBFF_SUPPORT (PF0_DEV_CAP2_OBFF_SUPPORT),
    .PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT (PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT),
    .PF0_DEV_CAP_ENDPOINT_L0S_LATENCY (PF0_DEV_CAP_ENDPOINT_L0S_LATENCY),
    .PF0_DEV_CAP_ENDPOINT_L1_LATENCY (PF0_DEV_CAP_ENDPOINT_L1_LATENCY),
    .PF0_DEV_CAP_EXT_TAG_SUPPORTED (PF0_DEV_CAP_EXT_TAG_SUPPORTED),
    .PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE (PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE),
    .PF0_DEV_CAP_MAX_PAYLOAD_SIZE (PF0_DEV_CAP_MAX_PAYLOAD_SIZE),
    .PF0_DPA_CAP_NEXTPTR (PF0_DPA_CAP_NEXTPTR),
    .PF0_DPA_CAP_SUB_STATE_CONTROL (PF0_DPA_CAP_SUB_STATE_CONTROL),
    .PF0_DPA_CAP_SUB_STATE_CONTROL_EN (PF0_DPA_CAP_SUB_STATE_CONTROL_EN),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6),
    .PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 (PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7),
    .PF0_DPA_CAP_VER (PF0_DPA_CAP_VER),
    .PF0_DSN_CAP_NEXTPTR (PF0_DSN_CAP_NEXTPTR),
    .PF0_EXPANSION_ROM_APERTURE_SIZE (PF0_EXPANSION_ROM_APERTURE_SIZE),
    .PF0_EXPANSION_ROM_ENABLE (PF0_EXPANSION_ROM_ENABLE),
    .PF0_INTERRUPT_LINE (PF0_INTERRUPT_LINE),
    .PF0_INTERRUPT_PIN (PF0_INTERRUPT_PIN),
    .PF0_LINK_CAP_ASPM_SUPPORT (PF0_LINK_CAP_ASPM_SUPPORT),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 (PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2),
    .PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 (PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 (PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2),
    .PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 (PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3),
    .PF0_LINK_STATUS_SLOT_CLOCK_CONFIG (PF0_LINK_STATUS_SLOT_CLOCK_CONFIG),
    .PF0_LTR_CAP_MAX_NOSNOOP_LAT (PF0_LTR_CAP_MAX_NOSNOOP_LAT),
    .PF0_LTR_CAP_MAX_SNOOP_LAT (PF0_LTR_CAP_MAX_SNOOP_LAT),
    .PF0_LTR_CAP_NEXTPTR (PF0_LTR_CAP_NEXTPTR),
    .PF0_LTR_CAP_VER (PF0_LTR_CAP_VER),
    .PF0_MSIX_CAP_NEXTPTR (PF0_MSIX_CAP_NEXTPTR),
    .PF0_MSIX_CAP_PBA_BIR (PF0_MSIX_CAP_PBA_BIR),
    .PF0_MSIX_CAP_PBA_OFFSET (PF0_MSIX_CAP_PBA_OFFSET),
    .PF0_MSIX_CAP_TABLE_BIR (PF0_MSIX_CAP_TABLE_BIR),
    .PF0_MSIX_CAP_TABLE_OFFSET (PF0_MSIX_CAP_TABLE_OFFSET),
    .PF0_MSIX_CAP_TABLE_SIZE (PF0_MSIX_CAP_TABLE_SIZE),
    .PF0_MSI_CAP_MULTIMSGCAP (PF0_MSI_CAP_MULTIMSGCAP),
    .PF0_MSI_CAP_NEXTPTR (PF0_MSI_CAP_NEXTPTR),
    .PF0_PB_CAP_NEXTPTR (PF0_PB_CAP_NEXTPTR),
    .PF0_PB_CAP_SYSTEM_ALLOCATED (PF0_PB_CAP_SYSTEM_ALLOCATED),
    .PF0_PB_CAP_VER (PF0_PB_CAP_VER),
    .PF0_PM_CAP_ID (PF0_PM_CAP_ID),
    .PF0_PM_CAP_NEXTPTR (PF0_PM_CAP_NEXTPTR),
    .PF0_PM_CAP_PMESUPPORT_D0 (PF0_PM_CAP_PMESUPPORT_D0),
    .PF0_PM_CAP_PMESUPPORT_D1 (PF0_PM_CAP_PMESUPPORT_D1),
    .PF0_PM_CAP_PMESUPPORT_D3HOT (PF0_PM_CAP_PMESUPPORT_D3HOT),
    .PF0_PM_CAP_SUPP_D1_STATE (PF0_PM_CAP_SUPP_D1_STATE),
    .PF0_PM_CAP_VER_ID (PF0_PM_CAP_VER_ID),
    .PF0_PM_CSR_NOSOFTRESET (PF0_PM_CSR_NOSOFTRESET),
    .PF0_RBAR_CAP_ENABLE (PF0_RBAR_CAP_ENABLE),
    .PF0_RBAR_CAP_INDEX0 (PF0_RBAR_CAP_INDEX0),
    .PF0_RBAR_CAP_INDEX1 (PF0_RBAR_CAP_INDEX1),
    .PF0_RBAR_CAP_INDEX2 (PF0_RBAR_CAP_INDEX2),
    .PF0_RBAR_CAP_NEXTPTR (PF0_RBAR_CAP_NEXTPTR),
    .PF0_RBAR_CAP_SIZE0 (PF0_RBAR_CAP_SIZE0),
    .PF0_RBAR_CAP_SIZE1 (PF0_RBAR_CAP_SIZE1),
    .PF0_RBAR_CAP_SIZE2 (PF0_RBAR_CAP_SIZE2),
    .PF0_RBAR_CAP_VER (PF0_RBAR_CAP_VER),
    .PF0_RBAR_NUM (PF0_RBAR_NUM),
    .PF0_REVISION_ID (PF0_REVISION_ID),
    .PF0_SRIOV_BAR0_APERTURE_SIZE (PF0_SRIOV_BAR0_APERTURE_SIZE),
    .PF0_SRIOV_BAR0_CONTROL (PF0_SRIOV_BAR0_CONTROL),
    .PF0_SRIOV_BAR1_APERTURE_SIZE (PF0_SRIOV_BAR1_APERTURE_SIZE),
    .PF0_SRIOV_BAR1_CONTROL (PF0_SRIOV_BAR1_CONTROL),
    .PF0_SRIOV_BAR2_APERTURE_SIZE (PF0_SRIOV_BAR2_APERTURE_SIZE),
    .PF0_SRIOV_BAR2_CONTROL (PF0_SRIOV_BAR2_CONTROL),
    .PF0_SRIOV_BAR3_APERTURE_SIZE (PF0_SRIOV_BAR3_APERTURE_SIZE),
    .PF0_SRIOV_BAR3_CONTROL (PF0_SRIOV_BAR3_CONTROL),
    .PF0_SRIOV_BAR4_APERTURE_SIZE (PF0_SRIOV_BAR4_APERTURE_SIZE),
    .PF0_SRIOV_BAR4_CONTROL (PF0_SRIOV_BAR4_CONTROL),
    .PF0_SRIOV_BAR5_APERTURE_SIZE (PF0_SRIOV_BAR5_APERTURE_SIZE),
    .PF0_SRIOV_BAR5_CONTROL (PF0_SRIOV_BAR5_CONTROL),
    .PF0_SRIOV_CAP_INITIAL_VF (PF0_SRIOV_CAP_INITIAL_VF),
    .PF0_SRIOV_CAP_NEXTPTR (PF0_SRIOV_CAP_NEXTPTR),
    .PF0_SRIOV_CAP_TOTAL_VF (PF0_SRIOV_CAP_TOTAL_VF),
    .PF0_SRIOV_CAP_VER (PF0_SRIOV_CAP_VER),
    .PF0_SRIOV_FIRST_VF_OFFSET (PF0_SRIOV_FIRST_VF_OFFSET),
    .PF0_SRIOV_FUNC_DEP_LINK (PF0_SRIOV_FUNC_DEP_LINK),
    .PF0_SRIOV_SUPPORTED_PAGE_SIZE (PF0_SRIOV_SUPPORTED_PAGE_SIZE),
    .PF0_SRIOV_VF_DEVICE_ID (PF0_SRIOV_VF_DEVICE_ID),
    .PF0_SUBSYSTEM_ID (PF0_SUBSYSTEM_ID),
    .PF0_TPHR_CAP_DEV_SPECIFIC_MODE (PF0_TPHR_CAP_DEV_SPECIFIC_MODE),
    .PF0_TPHR_CAP_ENABLE (PF0_TPHR_CAP_ENABLE),
    .PF0_TPHR_CAP_INT_VEC_MODE (PF0_TPHR_CAP_INT_VEC_MODE),
    .PF0_TPHR_CAP_NEXTPTR (PF0_TPHR_CAP_NEXTPTR),
    .PF0_TPHR_CAP_ST_MODE_SEL (PF0_TPHR_CAP_ST_MODE_SEL),
    .PF0_TPHR_CAP_ST_TABLE_LOC (PF0_TPHR_CAP_ST_TABLE_LOC),
    .PF0_TPHR_CAP_ST_TABLE_SIZE (PF0_TPHR_CAP_ST_TABLE_SIZE),
    .PF0_TPHR_CAP_VER (PF0_TPHR_CAP_VER),
    .PF0_VC_CAP_NEXTPTR (PF0_VC_CAP_NEXTPTR),
    .PF0_VC_CAP_VER (PF0_VC_CAP_VER),
    .PF1_AER_CAP_ECRC_CHECK_CAPABLE (PF1_AER_CAP_ECRC_CHECK_CAPABLE),
    .PF1_AER_CAP_ECRC_GEN_CAPABLE (PF1_AER_CAP_ECRC_GEN_CAPABLE),
    .PF1_AER_CAP_NEXTPTR (PF1_AER_CAP_NEXTPTR),
    .PF1_ARI_CAP_NEXTPTR (PF1_ARI_CAP_NEXTPTR),
    .PF1_ARI_CAP_NEXT_FUNC (PF1_ARI_CAP_NEXT_FUNC),
    .PF1_BAR0_APERTURE_SIZE (PF1_BAR0_APERTURE_SIZE),
    .PF1_BAR0_CONTROL (PF1_BAR0_CONTROL),
    .PF1_BAR1_APERTURE_SIZE (PF1_BAR1_APERTURE_SIZE),
    .PF1_BAR1_CONTROL (PF1_BAR1_CONTROL),
    .PF1_BAR2_APERTURE_SIZE (PF1_BAR2_APERTURE_SIZE),
    .PF1_BAR2_CONTROL (PF1_BAR2_CONTROL),
    .PF1_BAR3_APERTURE_SIZE (PF1_BAR3_APERTURE_SIZE),
    .PF1_BAR3_CONTROL (PF1_BAR3_CONTROL),
    .PF1_BAR4_APERTURE_SIZE (PF1_BAR4_APERTURE_SIZE),
    .PF1_BAR4_CONTROL (PF1_BAR4_CONTROL),
    .PF1_BAR5_APERTURE_SIZE (PF1_BAR5_APERTURE_SIZE),
    .PF1_BAR5_CONTROL (PF1_BAR5_CONTROL),
    .PF1_BIST_REGISTER (PF1_BIST_REGISTER),
    .PF1_CAPABILITY_POINTER (PF1_CAPABILITY_POINTER),
    .PF1_CLASS_CODE (PF1_CLASS_CODE),
    .PF1_DEVICE_ID (PF1_DEVICE_ID),
    .PF1_DEV_CAP_MAX_PAYLOAD_SIZE (PF1_DEV_CAP_MAX_PAYLOAD_SIZE),
    .PF1_DPA_CAP_NEXTPTR (PF1_DPA_CAP_NEXTPTR),
    .PF1_DPA_CAP_SUB_STATE_CONTROL (PF1_DPA_CAP_SUB_STATE_CONTROL),
    .PF1_DPA_CAP_SUB_STATE_CONTROL_EN (PF1_DPA_CAP_SUB_STATE_CONTROL_EN),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6),
    .PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 (PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7),
    .PF1_DPA_CAP_VER (PF1_DPA_CAP_VER),
    .PF1_DSN_CAP_NEXTPTR (PF1_DSN_CAP_NEXTPTR),
    .PF1_EXPANSION_ROM_APERTURE_SIZE (PF1_EXPANSION_ROM_APERTURE_SIZE),
    .PF1_EXPANSION_ROM_ENABLE (PF1_EXPANSION_ROM_ENABLE),
    .PF1_INTERRUPT_LINE (PF1_INTERRUPT_LINE),
    .PF1_INTERRUPT_PIN (PF1_INTERRUPT_PIN),
    .PF1_MSIX_CAP_NEXTPTR (PF1_MSIX_CAP_NEXTPTR),
    .PF1_MSIX_CAP_PBA_BIR (PF1_MSIX_CAP_PBA_BIR),
    .PF1_MSIX_CAP_PBA_OFFSET (PF1_MSIX_CAP_PBA_OFFSET),
    .PF1_MSIX_CAP_TABLE_BIR (PF1_MSIX_CAP_TABLE_BIR),
    .PF1_MSIX_CAP_TABLE_OFFSET (PF1_MSIX_CAP_TABLE_OFFSET),
    .PF1_MSIX_CAP_TABLE_SIZE (PF1_MSIX_CAP_TABLE_SIZE),
    .PF1_MSI_CAP_MULTIMSGCAP (PF1_MSI_CAP_MULTIMSGCAP),
    .PF1_MSI_CAP_NEXTPTR (PF1_MSI_CAP_NEXTPTR),
    .PF1_PB_CAP_NEXTPTR (PF1_PB_CAP_NEXTPTR),
    .PF1_PB_CAP_SYSTEM_ALLOCATED (PF1_PB_CAP_SYSTEM_ALLOCATED),
    .PF1_PB_CAP_VER (PF1_PB_CAP_VER),
    .PF1_PM_CAP_ID (PF1_PM_CAP_ID),
    .PF1_PM_CAP_NEXTPTR (PF1_PM_CAP_NEXTPTR),
    .PF1_PM_CAP_VER_ID (PF1_PM_CAP_VER_ID),
    .PF1_RBAR_CAP_ENABLE (PF1_RBAR_CAP_ENABLE),
    .PF1_RBAR_CAP_INDEX0 (PF1_RBAR_CAP_INDEX0),
    .PF1_RBAR_CAP_INDEX1 (PF1_RBAR_CAP_INDEX1),
    .PF1_RBAR_CAP_INDEX2 (PF1_RBAR_CAP_INDEX2),
    .PF1_RBAR_CAP_NEXTPTR (PF1_RBAR_CAP_NEXTPTR),
    .PF1_RBAR_CAP_SIZE0 (PF1_RBAR_CAP_SIZE0),
    .PF1_RBAR_CAP_SIZE1 (PF1_RBAR_CAP_SIZE1),
    .PF1_RBAR_CAP_SIZE2 (PF1_RBAR_CAP_SIZE2),
    .PF1_RBAR_CAP_VER (PF1_RBAR_CAP_VER),
    .PF1_RBAR_NUM (PF1_RBAR_NUM),
    .PF1_REVISION_ID (PF1_REVISION_ID),
    .PF1_SRIOV_BAR0_APERTURE_SIZE (PF1_SRIOV_BAR0_APERTURE_SIZE),
    .PF1_SRIOV_BAR0_CONTROL (PF1_SRIOV_BAR0_CONTROL),
    .PF1_SRIOV_BAR1_APERTURE_SIZE (PF1_SRIOV_BAR1_APERTURE_SIZE),
    .PF1_SRIOV_BAR1_CONTROL (PF1_SRIOV_BAR1_CONTROL),
    .PF1_SRIOV_BAR2_APERTURE_SIZE (PF1_SRIOV_BAR2_APERTURE_SIZE),
    .PF1_SRIOV_BAR2_CONTROL (PF1_SRIOV_BAR2_CONTROL),
    .PF1_SRIOV_BAR3_APERTURE_SIZE (PF1_SRIOV_BAR3_APERTURE_SIZE),
    .PF1_SRIOV_BAR3_CONTROL (PF1_SRIOV_BAR3_CONTROL),
    .PF1_SRIOV_BAR4_APERTURE_SIZE (PF1_SRIOV_BAR4_APERTURE_SIZE),
    .PF1_SRIOV_BAR4_CONTROL (PF1_SRIOV_BAR4_CONTROL),
    .PF1_SRIOV_BAR5_APERTURE_SIZE (PF1_SRIOV_BAR5_APERTURE_SIZE),
    .PF1_SRIOV_BAR5_CONTROL (PF1_SRIOV_BAR5_CONTROL),
    .PF1_SRIOV_CAP_INITIAL_VF (PF1_SRIOV_CAP_INITIAL_VF),
    .PF1_SRIOV_CAP_NEXTPTR (PF1_SRIOV_CAP_NEXTPTR),
    .PF1_SRIOV_CAP_TOTAL_VF (PF1_SRIOV_CAP_TOTAL_VF),
    .PF1_SRIOV_CAP_VER (PF1_SRIOV_CAP_VER),
    .PF1_SRIOV_FIRST_VF_OFFSET (PF1_SRIOV_FIRST_VF_OFFSET),
    .PF1_SRIOV_FUNC_DEP_LINK (PF1_SRIOV_FUNC_DEP_LINK),
    .PF1_SRIOV_SUPPORTED_PAGE_SIZE (PF1_SRIOV_SUPPORTED_PAGE_SIZE),
    .PF1_SRIOV_VF_DEVICE_ID (PF1_SRIOV_VF_DEVICE_ID),
    .PF1_SUBSYSTEM_ID (PF1_SUBSYSTEM_ID),
    .PF1_TPHR_CAP_DEV_SPECIFIC_MODE (PF1_TPHR_CAP_DEV_SPECIFIC_MODE),
    .PF1_TPHR_CAP_ENABLE (PF1_TPHR_CAP_ENABLE),
    .PF1_TPHR_CAP_INT_VEC_MODE (PF1_TPHR_CAP_INT_VEC_MODE),
    .PF1_TPHR_CAP_NEXTPTR (PF1_TPHR_CAP_NEXTPTR),
    .PF1_TPHR_CAP_ST_MODE_SEL (PF1_TPHR_CAP_ST_MODE_SEL),
    .PF1_TPHR_CAP_ST_TABLE_LOC (PF1_TPHR_CAP_ST_TABLE_LOC),
    .PF1_TPHR_CAP_ST_TABLE_SIZE (PF1_TPHR_CAP_ST_TABLE_SIZE),
    .PF1_TPHR_CAP_VER (PF1_TPHR_CAP_VER),
    .PL_DISABLE_EI_INFER_IN_L0 (PL_DISABLE_EI_INFER_IN_L0),
    .PL_DISABLE_GEN3_DC_BALANCE (PL_DISABLE_GEN3_DC_BALANCE),
    .PL_DISABLE_SCRAMBLING (PL_DISABLE_SCRAMBLING),
    .PL_DISABLE_UPCONFIG_CAPABLE (PL_DISABLE_UPCONFIG_CAPABLE),
    .PL_EQ_ADAPT_DISABLE_COEFF_CHECK (PL_EQ_ADAPT_DISABLE_COEFF_CHECK),
    .PL_EQ_ADAPT_DISABLE_PRESET_CHECK (PL_EQ_ADAPT_DISABLE_PRESET_CHECK),
    .PL_EQ_ADAPT_ITER_COUNT (PL_EQ_ADAPT_ITER_COUNT),
    .PL_EQ_ADAPT_REJECT_RETRY_COUNT (PL_EQ_ADAPT_REJECT_RETRY_COUNT),
    .PL_EQ_BYPASS_PHASE23 (PL_EQ_BYPASS_PHASE23),
    .PL_EQ_SHORT_ADAPT_PHASE (PL_EQ_SHORT_ADAPT_PHASE),
    .PL_LANE0_EQ_CONTROL (PL_LANE0_EQ_CONTROL),
    .PL_LANE1_EQ_CONTROL (PL_LANE1_EQ_CONTROL),
    .PL_LANE2_EQ_CONTROL (PL_LANE2_EQ_CONTROL),
    .PL_LANE3_EQ_CONTROL (PL_LANE3_EQ_CONTROL),
    .PL_LANE4_EQ_CONTROL (PL_LANE4_EQ_CONTROL),
    .PL_LANE5_EQ_CONTROL (PL_LANE5_EQ_CONTROL),
    .PL_LANE6_EQ_CONTROL (PL_LANE6_EQ_CONTROL),
    .PL_LANE7_EQ_CONTROL (PL_LANE7_EQ_CONTROL),
    .PL_LINK_CAP_MAX_LINK_SPEED (PL_LINK_CAP_MAX_LINK_SPEED),
    .PL_LINK_CAP_MAX_LINK_WIDTH (PL_LINK_CAP_MAX_LINK_WIDTH),
    .PL_N_FTS_COMCLK_GEN1 (PL_N_FTS_COMCLK_GEN1),
    .PL_N_FTS_COMCLK_GEN2 (PL_N_FTS_COMCLK_GEN2),
    .PL_N_FTS_COMCLK_GEN3 (PL_N_FTS_COMCLK_GEN3),
    .PL_N_FTS_GEN1 (PL_N_FTS_GEN1),
    .PL_N_FTS_GEN2 (PL_N_FTS_GEN2),
    .PL_N_FTS_GEN3 (PL_N_FTS_GEN3),
    .PL_SIM_FAST_LINK_TRAINING (PL_SIM_FAST_LINK_TRAINING),
    .PL_UPSTREAM_FACING (PL_UPSTREAM_FACING),
    .PM_ASPML0S_TIMEOUT (PM_ASPML0S_TIMEOUT),
    .PM_ASPML1_ENTRY_DELAY (PM_ASPML1_ENTRY_DELAY),
    .PM_ENABLE_SLOT_POWER_CAPTURE (PM_ENABLE_SLOT_POWER_CAPTURE),
    .PM_L1_REENTRY_DELAY (PM_L1_REENTRY_DELAY),
    .PM_PME_SERVICE_TIMEOUT_DELAY (PM_PME_SERVICE_TIMEOUT_DELAY),
    .PM_PME_TURNOFF_ACK_DELAY (PM_PME_TURNOFF_ACK_DELAY),
    .SIM_VERSION (SIM_VERSION),
    .SPARE_BIT0 (SPARE_BIT0),
    .SPARE_BIT1 (SPARE_BIT1),
    .SPARE_BIT2 (SPARE_BIT2),
    .SPARE_BIT3 (SPARE_BIT3),
    .SPARE_BIT4 (SPARE_BIT4),
    .SPARE_BIT5 (SPARE_BIT5),
    .SPARE_BIT6 (SPARE_BIT6),
    .SPARE_BIT7 (SPARE_BIT7),
    .SPARE_BIT8 (SPARE_BIT8),
    .SPARE_BYTE0 (SPARE_BYTE0),
    .SPARE_BYTE1 (SPARE_BYTE1),
    .SPARE_BYTE2 (SPARE_BYTE2),
    .SPARE_BYTE3 (SPARE_BYTE3),
    .SPARE_WORD0 (SPARE_WORD0),
    .SPARE_WORD1 (SPARE_WORD1),
    .SPARE_WORD2 (SPARE_WORD2),
    .SPARE_WORD3 (SPARE_WORD3),
    .SRIOV_CAP_ENABLE (SRIOV_CAP_ENABLE),
    .TL_COMPL_TIMEOUT_REG0 (TL_COMPL_TIMEOUT_REG0),
    .TL_COMPL_TIMEOUT_REG1 (TL_COMPL_TIMEOUT_REG1),
    .TL_CREDITS_CD (TL_CREDITS_CD),
    .TL_CREDITS_CH (TL_CREDITS_CH),
    .TL_CREDITS_NPD (TL_CREDITS_NPD),
    .TL_CREDITS_NPH (TL_CREDITS_NPH),
    .TL_CREDITS_PD (TL_CREDITS_PD),
    .TL_CREDITS_PH (TL_CREDITS_PH),
    .TL_ENABLE_MESSAGE_RID_CHECK_ENABLE (TL_ENABLE_MESSAGE_RID_CHECK_ENABLE),
    .TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE (TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE),
    .TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE (TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE),
    .TL_LEGACY_MODE_ENABLE (TL_LEGACY_MODE_ENABLE),
    .TL_PF_ENABLE_REG (TL_PF_ENABLE_REG),
    .TL_TAG_MGMT_ENABLE (TL_TAG_MGMT_ENABLE),
    .VF0_ARI_CAP_NEXTPTR (VF0_ARI_CAP_NEXTPTR),
    .VF0_CAPABILITY_POINTER (VF0_CAPABILITY_POINTER),
    .VF0_MSIX_CAP_PBA_BIR (VF0_MSIX_CAP_PBA_BIR),
    .VF0_MSIX_CAP_PBA_OFFSET (VF0_MSIX_CAP_PBA_OFFSET),
    .VF0_MSIX_CAP_TABLE_BIR (VF0_MSIX_CAP_TABLE_BIR),
    .VF0_MSIX_CAP_TABLE_OFFSET (VF0_MSIX_CAP_TABLE_OFFSET),
    .VF0_MSIX_CAP_TABLE_SIZE (VF0_MSIX_CAP_TABLE_SIZE),
    .VF0_MSI_CAP_MULTIMSGCAP (VF0_MSI_CAP_MULTIMSGCAP),
    .VF0_PM_CAP_ID (VF0_PM_CAP_ID),
    .VF0_PM_CAP_NEXTPTR (VF0_PM_CAP_NEXTPTR),
    .VF0_PM_CAP_VER_ID (VF0_PM_CAP_VER_ID),
    .VF0_TPHR_CAP_DEV_SPECIFIC_MODE (VF0_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF0_TPHR_CAP_ENABLE (VF0_TPHR_CAP_ENABLE),
    .VF0_TPHR_CAP_INT_VEC_MODE (VF0_TPHR_CAP_INT_VEC_MODE),
    .VF0_TPHR_CAP_NEXTPTR (VF0_TPHR_CAP_NEXTPTR),
    .VF0_TPHR_CAP_ST_MODE_SEL (VF0_TPHR_CAP_ST_MODE_SEL),
    .VF0_TPHR_CAP_ST_TABLE_LOC (VF0_TPHR_CAP_ST_TABLE_LOC),
    .VF0_TPHR_CAP_ST_TABLE_SIZE (VF0_TPHR_CAP_ST_TABLE_SIZE),
    .VF0_TPHR_CAP_VER (VF0_TPHR_CAP_VER),
    .VF1_ARI_CAP_NEXTPTR (VF1_ARI_CAP_NEXTPTR),
    .VF1_MSIX_CAP_PBA_BIR (VF1_MSIX_CAP_PBA_BIR),
    .VF1_MSIX_CAP_PBA_OFFSET (VF1_MSIX_CAP_PBA_OFFSET),
    .VF1_MSIX_CAP_TABLE_BIR (VF1_MSIX_CAP_TABLE_BIR),
    .VF1_MSIX_CAP_TABLE_OFFSET (VF1_MSIX_CAP_TABLE_OFFSET),
    .VF1_MSIX_CAP_TABLE_SIZE (VF1_MSIX_CAP_TABLE_SIZE),
    .VF1_MSI_CAP_MULTIMSGCAP (VF1_MSI_CAP_MULTIMSGCAP),
    .VF1_PM_CAP_ID (VF1_PM_CAP_ID),
    .VF1_PM_CAP_NEXTPTR (VF1_PM_CAP_NEXTPTR),
    .VF1_PM_CAP_VER_ID (VF1_PM_CAP_VER_ID),
    .VF1_TPHR_CAP_DEV_SPECIFIC_MODE (VF1_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF1_TPHR_CAP_ENABLE (VF1_TPHR_CAP_ENABLE),
    .VF1_TPHR_CAP_INT_VEC_MODE (VF1_TPHR_CAP_INT_VEC_MODE),
    .VF1_TPHR_CAP_NEXTPTR (VF1_TPHR_CAP_NEXTPTR),
    .VF1_TPHR_CAP_ST_MODE_SEL (VF1_TPHR_CAP_ST_MODE_SEL),
    .VF1_TPHR_CAP_ST_TABLE_LOC (VF1_TPHR_CAP_ST_TABLE_LOC),
    .VF1_TPHR_CAP_ST_TABLE_SIZE (VF1_TPHR_CAP_ST_TABLE_SIZE),
    .VF1_TPHR_CAP_VER (VF1_TPHR_CAP_VER),
    .VF2_ARI_CAP_NEXTPTR (VF2_ARI_CAP_NEXTPTR),
    .VF2_MSIX_CAP_PBA_BIR (VF2_MSIX_CAP_PBA_BIR),
    .VF2_MSIX_CAP_PBA_OFFSET (VF2_MSIX_CAP_PBA_OFFSET),
    .VF2_MSIX_CAP_TABLE_BIR (VF2_MSIX_CAP_TABLE_BIR),
    .VF2_MSIX_CAP_TABLE_OFFSET (VF2_MSIX_CAP_TABLE_OFFSET),
    .VF2_MSIX_CAP_TABLE_SIZE (VF2_MSIX_CAP_TABLE_SIZE),
    .VF2_MSI_CAP_MULTIMSGCAP (VF2_MSI_CAP_MULTIMSGCAP),
    .VF2_PM_CAP_ID (VF2_PM_CAP_ID),
    .VF2_PM_CAP_NEXTPTR (VF2_PM_CAP_NEXTPTR),
    .VF2_PM_CAP_VER_ID (VF2_PM_CAP_VER_ID),
    .VF2_TPHR_CAP_DEV_SPECIFIC_MODE (VF2_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF2_TPHR_CAP_ENABLE (VF2_TPHR_CAP_ENABLE),
    .VF2_TPHR_CAP_INT_VEC_MODE (VF2_TPHR_CAP_INT_VEC_MODE),
    .VF2_TPHR_CAP_NEXTPTR (VF2_TPHR_CAP_NEXTPTR),
    .VF2_TPHR_CAP_ST_MODE_SEL (VF2_TPHR_CAP_ST_MODE_SEL),
    .VF2_TPHR_CAP_ST_TABLE_LOC (VF2_TPHR_CAP_ST_TABLE_LOC),
    .VF2_TPHR_CAP_ST_TABLE_SIZE (VF2_TPHR_CAP_ST_TABLE_SIZE),
    .VF2_TPHR_CAP_VER (VF2_TPHR_CAP_VER),
    .VF3_ARI_CAP_NEXTPTR (VF3_ARI_CAP_NEXTPTR),
    .VF3_MSIX_CAP_PBA_BIR (VF3_MSIX_CAP_PBA_BIR),
    .VF3_MSIX_CAP_PBA_OFFSET (VF3_MSIX_CAP_PBA_OFFSET),
    .VF3_MSIX_CAP_TABLE_BIR (VF3_MSIX_CAP_TABLE_BIR),
    .VF3_MSIX_CAP_TABLE_OFFSET (VF3_MSIX_CAP_TABLE_OFFSET),
    .VF3_MSIX_CAP_TABLE_SIZE (VF3_MSIX_CAP_TABLE_SIZE),
    .VF3_MSI_CAP_MULTIMSGCAP (VF3_MSI_CAP_MULTIMSGCAP),
    .VF3_PM_CAP_ID (VF3_PM_CAP_ID),
    .VF3_PM_CAP_NEXTPTR (VF3_PM_CAP_NEXTPTR),
    .VF3_PM_CAP_VER_ID (VF3_PM_CAP_VER_ID),
    .VF3_TPHR_CAP_DEV_SPECIFIC_MODE (VF3_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF3_TPHR_CAP_ENABLE (VF3_TPHR_CAP_ENABLE),
    .VF3_TPHR_CAP_INT_VEC_MODE (VF3_TPHR_CAP_INT_VEC_MODE),
    .VF3_TPHR_CAP_NEXTPTR (VF3_TPHR_CAP_NEXTPTR),
    .VF3_TPHR_CAP_ST_MODE_SEL (VF3_TPHR_CAP_ST_MODE_SEL),
    .VF3_TPHR_CAP_ST_TABLE_LOC (VF3_TPHR_CAP_ST_TABLE_LOC),
    .VF3_TPHR_CAP_ST_TABLE_SIZE (VF3_TPHR_CAP_ST_TABLE_SIZE),
    .VF3_TPHR_CAP_VER (VF3_TPHR_CAP_VER),
    .VF4_ARI_CAP_NEXTPTR (VF4_ARI_CAP_NEXTPTR),
    .VF4_MSIX_CAP_PBA_BIR (VF4_MSIX_CAP_PBA_BIR),
    .VF4_MSIX_CAP_PBA_OFFSET (VF4_MSIX_CAP_PBA_OFFSET),
    .VF4_MSIX_CAP_TABLE_BIR (VF4_MSIX_CAP_TABLE_BIR),
    .VF4_MSIX_CAP_TABLE_OFFSET (VF4_MSIX_CAP_TABLE_OFFSET),
    .VF4_MSIX_CAP_TABLE_SIZE (VF4_MSIX_CAP_TABLE_SIZE),
    .VF4_MSI_CAP_MULTIMSGCAP (VF4_MSI_CAP_MULTIMSGCAP),
    .VF4_PM_CAP_ID (VF4_PM_CAP_ID),
    .VF4_PM_CAP_NEXTPTR (VF4_PM_CAP_NEXTPTR),
    .VF4_PM_CAP_VER_ID (VF4_PM_CAP_VER_ID),
    .VF4_TPHR_CAP_DEV_SPECIFIC_MODE (VF4_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF4_TPHR_CAP_ENABLE (VF4_TPHR_CAP_ENABLE),
    .VF4_TPHR_CAP_INT_VEC_MODE (VF4_TPHR_CAP_INT_VEC_MODE),
    .VF4_TPHR_CAP_NEXTPTR (VF4_TPHR_CAP_NEXTPTR),
    .VF4_TPHR_CAP_ST_MODE_SEL (VF4_TPHR_CAP_ST_MODE_SEL),
    .VF4_TPHR_CAP_ST_TABLE_LOC (VF4_TPHR_CAP_ST_TABLE_LOC),
    .VF4_TPHR_CAP_ST_TABLE_SIZE (VF4_TPHR_CAP_ST_TABLE_SIZE),
    .VF4_TPHR_CAP_VER (VF4_TPHR_CAP_VER),
    .VF5_ARI_CAP_NEXTPTR (VF5_ARI_CAP_NEXTPTR),
    .VF5_MSIX_CAP_PBA_BIR (VF5_MSIX_CAP_PBA_BIR),
    .VF5_MSIX_CAP_PBA_OFFSET (VF5_MSIX_CAP_PBA_OFFSET),
    .VF5_MSIX_CAP_TABLE_BIR (VF5_MSIX_CAP_TABLE_BIR),
    .VF5_MSIX_CAP_TABLE_OFFSET (VF5_MSIX_CAP_TABLE_OFFSET),
    .VF5_MSIX_CAP_TABLE_SIZE (VF5_MSIX_CAP_TABLE_SIZE),
    .VF5_MSI_CAP_MULTIMSGCAP (VF5_MSI_CAP_MULTIMSGCAP),
    .VF5_PM_CAP_ID (VF5_PM_CAP_ID),
    .VF5_PM_CAP_NEXTPTR (VF5_PM_CAP_NEXTPTR),
    .VF5_PM_CAP_VER_ID (VF5_PM_CAP_VER_ID),
    .VF5_TPHR_CAP_DEV_SPECIFIC_MODE (VF5_TPHR_CAP_DEV_SPECIFIC_MODE),
    .VF5_TPHR_CAP_ENABLE (VF5_TPHR_CAP_ENABLE),
    .VF5_TPHR_CAP_INT_VEC_MODE (VF5_TPHR_CAP_INT_VEC_MODE),
    .VF5_TPHR_CAP_NEXTPTR (VF5_TPHR_CAP_NEXTPTR),
    .VF5_TPHR_CAP_ST_MODE_SEL (VF5_TPHR_CAP_ST_MODE_SEL),
    .VF5_TPHR_CAP_ST_TABLE_LOC (VF5_TPHR_CAP_ST_TABLE_LOC),
    .VF5_TPHR_CAP_ST_TABLE_SIZE (VF5_TPHR_CAP_ST_TABLE_SIZE),
    .VF5_TPHR_CAP_VER (VF5_TPHR_CAP_VER))

    B_PCIE_3_0_INST (
    .CFGCURRENTSPEED (delay_CFGCURRENTSPEED),
    .CFGDPASUBSTATECHANGE (delay_CFGDPASUBSTATECHANGE),
    .CFGERRCOROUT (delay_CFGERRCOROUT),
    .CFGERRFATALOUT (delay_CFGERRFATALOUT),
    .CFGERRNONFATALOUT (delay_CFGERRNONFATALOUT),
    .CFGEXTFUNCTIONNUMBER (delay_CFGEXTFUNCTIONNUMBER),
    .CFGEXTREADRECEIVED (delay_CFGEXTREADRECEIVED),
    .CFGEXTREGISTERNUMBER (delay_CFGEXTREGISTERNUMBER),
    .CFGEXTWRITEBYTEENABLE (delay_CFGEXTWRITEBYTEENABLE),
    .CFGEXTWRITEDATA (delay_CFGEXTWRITEDATA),
    .CFGEXTWRITERECEIVED (delay_CFGEXTWRITERECEIVED),
    .CFGFCCPLD (delay_CFGFCCPLD),
    .CFGFCCPLH (delay_CFGFCCPLH),
    .CFGFCNPD (delay_CFGFCNPD),
    .CFGFCNPH (delay_CFGFCNPH),
    .CFGFCPD (delay_CFGFCPD),
    .CFGFCPH (delay_CFGFCPH),
    .CFGFLRINPROCESS (delay_CFGFLRINPROCESS),
    .CFGFUNCTIONPOWERSTATE (delay_CFGFUNCTIONPOWERSTATE),
    .CFGFUNCTIONSTATUS (delay_CFGFUNCTIONSTATUS),
    .CFGHOTRESETOUT (delay_CFGHOTRESETOUT),
    .CFGINPUTUPDATEDONE (delay_CFGINPUTUPDATEDONE),
    .CFGINTERRUPTAOUTPUT (delay_CFGINTERRUPTAOUTPUT),
    .CFGINTERRUPTBOUTPUT (delay_CFGINTERRUPTBOUTPUT),
    .CFGINTERRUPTCOUTPUT (delay_CFGINTERRUPTCOUTPUT),
    .CFGINTERRUPTDOUTPUT (delay_CFGINTERRUPTDOUTPUT),
    .CFGINTERRUPTMSIDATA (delay_CFGINTERRUPTMSIDATA),
    .CFGINTERRUPTMSIENABLE (delay_CFGINTERRUPTMSIENABLE),
    .CFGINTERRUPTMSIFAIL (delay_CFGINTERRUPTMSIFAIL),
    .CFGINTERRUPTMSIMASKUPDATE (delay_CFGINTERRUPTMSIMASKUPDATE),
    .CFGINTERRUPTMSIMMENABLE (delay_CFGINTERRUPTMSIMMENABLE),
    .CFGINTERRUPTMSISENT (delay_CFGINTERRUPTMSISENT),
    .CFGINTERRUPTMSIVFENABLE (delay_CFGINTERRUPTMSIVFENABLE),
    .CFGINTERRUPTMSIXENABLE (delay_CFGINTERRUPTMSIXENABLE),
    .CFGINTERRUPTMSIXFAIL (delay_CFGINTERRUPTMSIXFAIL),
    .CFGINTERRUPTMSIXMASK (delay_CFGINTERRUPTMSIXMASK),
    .CFGINTERRUPTMSIXSENT (delay_CFGINTERRUPTMSIXSENT),
    .CFGINTERRUPTMSIXVFENABLE (delay_CFGINTERRUPTMSIXVFENABLE),
    .CFGINTERRUPTMSIXVFMASK (delay_CFGINTERRUPTMSIXVFMASK),
    .CFGINTERRUPTSENT (delay_CFGINTERRUPTSENT),
    .CFGLINKPOWERSTATE (delay_CFGLINKPOWERSTATE),
    .CFGLOCALERROR (delay_CFGLOCALERROR),
    .CFGLTRENABLE (delay_CFGLTRENABLE),
    .CFGLTSSMSTATE (delay_CFGLTSSMSTATE),
    .CFGMAXPAYLOAD (delay_CFGMAXPAYLOAD),
    .CFGMAXREADREQ (delay_CFGMAXREADREQ),
    .CFGMCUPDATEDONE (delay_CFGMCUPDATEDONE),
    .CFGMGMTREADDATA (delay_CFGMGMTREADDATA),
    .CFGMGMTREADWRITEDONE (delay_CFGMGMTREADWRITEDONE),
    .CFGMSGRECEIVED (delay_CFGMSGRECEIVED),
    .CFGMSGRECEIVEDDATA (delay_CFGMSGRECEIVEDDATA),
    .CFGMSGRECEIVEDTYPE (delay_CFGMSGRECEIVEDTYPE),
    .CFGMSGTRANSMITDONE (delay_CFGMSGTRANSMITDONE),
    .CFGNEGOTIATEDWIDTH (delay_CFGNEGOTIATEDWIDTH),
    .CFGOBFFENABLE (delay_CFGOBFFENABLE),
    .CFGPERFUNCSTATUSDATA (delay_CFGPERFUNCSTATUSDATA),
    .CFGPERFUNCTIONUPDATEDONE (delay_CFGPERFUNCTIONUPDATEDONE),
    .CFGPHYLINKDOWN (delay_CFGPHYLINKDOWN),
    .CFGPHYLINKSTATUS (delay_CFGPHYLINKSTATUS),
    .CFGPLSTATUSCHANGE (delay_CFGPLSTATUSCHANGE),
    .CFGPOWERSTATECHANGEINTERRUPT (delay_CFGPOWERSTATECHANGEINTERRUPT),
    .CFGRCBSTATUS (delay_CFGRCBSTATUS),
    .CFGTPHFUNCTIONNUM (delay_CFGTPHFUNCTIONNUM),
    .CFGTPHREQUESTERENABLE (delay_CFGTPHREQUESTERENABLE),
    .CFGTPHSTMODE (delay_CFGTPHSTMODE),
    .CFGTPHSTTADDRESS (delay_CFGTPHSTTADDRESS),
    .CFGTPHSTTREADENABLE (delay_CFGTPHSTTREADENABLE),
    .CFGTPHSTTWRITEBYTEVALID (delay_CFGTPHSTTWRITEBYTEVALID),
    .CFGTPHSTTWRITEDATA (delay_CFGTPHSTTWRITEDATA),
    .CFGTPHSTTWRITEENABLE (delay_CFGTPHSTTWRITEENABLE),
    .CFGVFFLRINPROCESS (delay_CFGVFFLRINPROCESS),
    .CFGVFPOWERSTATE (delay_CFGVFPOWERSTATE),
    .CFGVFSTATUS (delay_CFGVFSTATUS),
    .CFGVFTPHREQUESTERENABLE (delay_CFGVFTPHREQUESTERENABLE),
    .CFGVFTPHSTMODE (delay_CFGVFTPHSTMODE),
    .DBGDATAOUT (delay_DBGDATAOUT),
    .DRPDO (delay_DRPDO),
    .DRPRDY (delay_DRPRDY),
    .MAXISCQTDATA (delay_MAXISCQTDATA),
    .MAXISCQTKEEP (delay_MAXISCQTKEEP),
    .MAXISCQTLAST (delay_MAXISCQTLAST),
    .MAXISCQTUSER (delay_MAXISCQTUSER),
    .MAXISCQTVALID (delay_MAXISCQTVALID),
    .MAXISRCTDATA (delay_MAXISRCTDATA),
    .MAXISRCTKEEP (delay_MAXISRCTKEEP),
    .MAXISRCTLAST (delay_MAXISRCTLAST),
    .MAXISRCTUSER (delay_MAXISRCTUSER),
    .MAXISRCTVALID (delay_MAXISRCTVALID),
    .MICOMPLETIONRAMREADADDRESSAL (delay_MICOMPLETIONRAMREADADDRESSAL),
    .MICOMPLETIONRAMREADADDRESSAU (delay_MICOMPLETIONRAMREADADDRESSAU),
    .MICOMPLETIONRAMREADADDRESSBL (delay_MICOMPLETIONRAMREADADDRESSBL),
    .MICOMPLETIONRAMREADADDRESSBU (delay_MICOMPLETIONRAMREADADDRESSBU),
    .MICOMPLETIONRAMREADENABLEL (delay_MICOMPLETIONRAMREADENABLEL),
    .MICOMPLETIONRAMREADENABLEU (delay_MICOMPLETIONRAMREADENABLEU),
    .MICOMPLETIONRAMWRITEADDRESSAL (delay_MICOMPLETIONRAMWRITEADDRESSAL),
    .MICOMPLETIONRAMWRITEADDRESSAU (delay_MICOMPLETIONRAMWRITEADDRESSAU),
    .MICOMPLETIONRAMWRITEADDRESSBL (delay_MICOMPLETIONRAMWRITEADDRESSBL),
    .MICOMPLETIONRAMWRITEADDRESSBU (delay_MICOMPLETIONRAMWRITEADDRESSBU),
    .MICOMPLETIONRAMWRITEDATAL (delay_MICOMPLETIONRAMWRITEDATAL),
    .MICOMPLETIONRAMWRITEDATAU (delay_MICOMPLETIONRAMWRITEDATAU),
    .MICOMPLETIONRAMWRITEENABLEL (delay_MICOMPLETIONRAMWRITEENABLEL),
    .MICOMPLETIONRAMWRITEENABLEU (delay_MICOMPLETIONRAMWRITEENABLEU),
    .MIREPLAYRAMADDRESS (delay_MIREPLAYRAMADDRESS),
    .MIREPLAYRAMREADENABLE (delay_MIREPLAYRAMREADENABLE),
    .MIREPLAYRAMWRITEDATA (delay_MIREPLAYRAMWRITEDATA),
    .MIREPLAYRAMWRITEENABLE (delay_MIREPLAYRAMWRITEENABLE),
    .MIREQUESTRAMREADADDRESSA (delay_MIREQUESTRAMREADADDRESSA),
    .MIREQUESTRAMREADADDRESSB (delay_MIREQUESTRAMREADADDRESSB),
    .MIREQUESTRAMREADENABLE (delay_MIREQUESTRAMREADENABLE),
    .MIREQUESTRAMWRITEADDRESSA (delay_MIREQUESTRAMWRITEADDRESSA),
    .MIREQUESTRAMWRITEADDRESSB (delay_MIREQUESTRAMWRITEADDRESSB),
    .MIREQUESTRAMWRITEDATA (delay_MIREQUESTRAMWRITEDATA),
    .MIREQUESTRAMWRITEENABLE (delay_MIREQUESTRAMWRITEENABLE),
    .PCIECQNPREQCOUNT (delay_PCIECQNPREQCOUNT),
    .PCIERQSEQNUM (delay_PCIERQSEQNUM),
    .PCIERQSEQNUMVLD (delay_PCIERQSEQNUMVLD),
    .PCIERQTAG (delay_PCIERQTAG),
    .PCIERQTAGAV (delay_PCIERQTAGAV),
    .PCIERQTAGVLD (delay_PCIERQTAGVLD),
    .PCIETFCNPDAV (delay_PCIETFCNPDAV),
    .PCIETFCNPHAV (delay_PCIETFCNPHAV),
    .PIPERX0EQCONTROL (delay_PIPERX0EQCONTROL),
    .PIPERX0EQLPLFFS (delay_PIPERX0EQLPLFFS),
    .PIPERX0EQLPTXPRESET (delay_PIPERX0EQLPTXPRESET),
    .PIPERX0EQPRESET (delay_PIPERX0EQPRESET),
    .PIPERX0POLARITY (delay_PIPERX0POLARITY),
    .PIPERX1EQCONTROL (delay_PIPERX1EQCONTROL),
    .PIPERX1EQLPLFFS (delay_PIPERX1EQLPLFFS),
    .PIPERX1EQLPTXPRESET (delay_PIPERX1EQLPTXPRESET),
    .PIPERX1EQPRESET (delay_PIPERX1EQPRESET),
    .PIPERX1POLARITY (delay_PIPERX1POLARITY),
    .PIPERX2EQCONTROL (delay_PIPERX2EQCONTROL),
    .PIPERX2EQLPLFFS (delay_PIPERX2EQLPLFFS),
    .PIPERX2EQLPTXPRESET (delay_PIPERX2EQLPTXPRESET),
    .PIPERX2EQPRESET (delay_PIPERX2EQPRESET),
    .PIPERX2POLARITY (delay_PIPERX2POLARITY),
    .PIPERX3EQCONTROL (delay_PIPERX3EQCONTROL),
    .PIPERX3EQLPLFFS (delay_PIPERX3EQLPLFFS),
    .PIPERX3EQLPTXPRESET (delay_PIPERX3EQLPTXPRESET),
    .PIPERX3EQPRESET (delay_PIPERX3EQPRESET),
    .PIPERX3POLARITY (delay_PIPERX3POLARITY),
    .PIPERX4EQCONTROL (delay_PIPERX4EQCONTROL),
    .PIPERX4EQLPLFFS (delay_PIPERX4EQLPLFFS),
    .PIPERX4EQLPTXPRESET (delay_PIPERX4EQLPTXPRESET),
    .PIPERX4EQPRESET (delay_PIPERX4EQPRESET),
    .PIPERX4POLARITY (delay_PIPERX4POLARITY),
    .PIPERX5EQCONTROL (delay_PIPERX5EQCONTROL),
    .PIPERX5EQLPLFFS (delay_PIPERX5EQLPLFFS),
    .PIPERX5EQLPTXPRESET (delay_PIPERX5EQLPTXPRESET),
    .PIPERX5EQPRESET (delay_PIPERX5EQPRESET),
    .PIPERX5POLARITY (delay_PIPERX5POLARITY),
    .PIPERX6EQCONTROL (delay_PIPERX6EQCONTROL),
    .PIPERX6EQLPLFFS (delay_PIPERX6EQLPLFFS),
    .PIPERX6EQLPTXPRESET (delay_PIPERX6EQLPTXPRESET),
    .PIPERX6EQPRESET (delay_PIPERX6EQPRESET),
    .PIPERX6POLARITY (delay_PIPERX6POLARITY),
    .PIPERX7EQCONTROL (delay_PIPERX7EQCONTROL),
    .PIPERX7EQLPLFFS (delay_PIPERX7EQLPLFFS),
    .PIPERX7EQLPTXPRESET (delay_PIPERX7EQLPTXPRESET),
    .PIPERX7EQPRESET (delay_PIPERX7EQPRESET),
    .PIPERX7POLARITY (delay_PIPERX7POLARITY),
    .PIPETX0CHARISK (delay_PIPETX0CHARISK),
    .PIPETX0COMPLIANCE (delay_PIPETX0COMPLIANCE),
    .PIPETX0DATA (delay_PIPETX0DATA),
    .PIPETX0DATAVALID (delay_PIPETX0DATAVALID),
    .PIPETX0ELECIDLE (delay_PIPETX0ELECIDLE),
    .PIPETX0EQCONTROL (delay_PIPETX0EQCONTROL),
    .PIPETX0EQDEEMPH (delay_PIPETX0EQDEEMPH),
    .PIPETX0EQPRESET (delay_PIPETX0EQPRESET),
    .PIPETX0POWERDOWN (delay_PIPETX0POWERDOWN),
    .PIPETX0STARTBLOCK (delay_PIPETX0STARTBLOCK),
    .PIPETX0SYNCHEADER (delay_PIPETX0SYNCHEADER),
    .PIPETX1CHARISK (delay_PIPETX1CHARISK),
    .PIPETX1COMPLIANCE (delay_PIPETX1COMPLIANCE),
    .PIPETX1DATA (delay_PIPETX1DATA),
    .PIPETX1DATAVALID (delay_PIPETX1DATAVALID),
    .PIPETX1ELECIDLE (delay_PIPETX1ELECIDLE),
    .PIPETX1EQCONTROL (delay_PIPETX1EQCONTROL),
    .PIPETX1EQDEEMPH (delay_PIPETX1EQDEEMPH),
    .PIPETX1EQPRESET (delay_PIPETX1EQPRESET),
    .PIPETX1POWERDOWN (delay_PIPETX1POWERDOWN),
    .PIPETX1STARTBLOCK (delay_PIPETX1STARTBLOCK),
    .PIPETX1SYNCHEADER (delay_PIPETX1SYNCHEADER),
    .PIPETX2CHARISK (delay_PIPETX2CHARISK),
    .PIPETX2COMPLIANCE (delay_PIPETX2COMPLIANCE),
    .PIPETX2DATA (delay_PIPETX2DATA),
    .PIPETX2DATAVALID (delay_PIPETX2DATAVALID),
    .PIPETX2ELECIDLE (delay_PIPETX2ELECIDLE),
    .PIPETX2EQCONTROL (delay_PIPETX2EQCONTROL),
    .PIPETX2EQDEEMPH (delay_PIPETX2EQDEEMPH),
    .PIPETX2EQPRESET (delay_PIPETX2EQPRESET),
    .PIPETX2POWERDOWN (delay_PIPETX2POWERDOWN),
    .PIPETX2STARTBLOCK (delay_PIPETX2STARTBLOCK),
    .PIPETX2SYNCHEADER (delay_PIPETX2SYNCHEADER),
    .PIPETX3CHARISK (delay_PIPETX3CHARISK),
    .PIPETX3COMPLIANCE (delay_PIPETX3COMPLIANCE),
    .PIPETX3DATA (delay_PIPETX3DATA),
    .PIPETX3DATAVALID (delay_PIPETX3DATAVALID),
    .PIPETX3ELECIDLE (delay_PIPETX3ELECIDLE),
    .PIPETX3EQCONTROL (delay_PIPETX3EQCONTROL),
    .PIPETX3EQDEEMPH (delay_PIPETX3EQDEEMPH),
    .PIPETX3EQPRESET (delay_PIPETX3EQPRESET),
    .PIPETX3POWERDOWN (delay_PIPETX3POWERDOWN),
    .PIPETX3STARTBLOCK (delay_PIPETX3STARTBLOCK),
    .PIPETX3SYNCHEADER (delay_PIPETX3SYNCHEADER),
    .PIPETX4CHARISK (delay_PIPETX4CHARISK),
    .PIPETX4COMPLIANCE (delay_PIPETX4COMPLIANCE),
    .PIPETX4DATA (delay_PIPETX4DATA),
    .PIPETX4DATAVALID (delay_PIPETX4DATAVALID),
    .PIPETX4ELECIDLE (delay_PIPETX4ELECIDLE),
    .PIPETX4EQCONTROL (delay_PIPETX4EQCONTROL),
    .PIPETX4EQDEEMPH (delay_PIPETX4EQDEEMPH),
    .PIPETX4EQPRESET (delay_PIPETX4EQPRESET),
    .PIPETX4POWERDOWN (delay_PIPETX4POWERDOWN),
    .PIPETX4STARTBLOCK (delay_PIPETX4STARTBLOCK),
    .PIPETX4SYNCHEADER (delay_PIPETX4SYNCHEADER),
    .PIPETX5CHARISK (delay_PIPETX5CHARISK),
    .PIPETX5COMPLIANCE (delay_PIPETX5COMPLIANCE),
    .PIPETX5DATA (delay_PIPETX5DATA),
    .PIPETX5DATAVALID (delay_PIPETX5DATAVALID),
    .PIPETX5ELECIDLE (delay_PIPETX5ELECIDLE),
    .PIPETX5EQCONTROL (delay_PIPETX5EQCONTROL),
    .PIPETX5EQDEEMPH (delay_PIPETX5EQDEEMPH),
    .PIPETX5EQPRESET (delay_PIPETX5EQPRESET),
    .PIPETX5POWERDOWN (delay_PIPETX5POWERDOWN),
    .PIPETX5STARTBLOCK (delay_PIPETX5STARTBLOCK),
    .PIPETX5SYNCHEADER (delay_PIPETX5SYNCHEADER),
    .PIPETX6CHARISK (delay_PIPETX6CHARISK),
    .PIPETX6COMPLIANCE (delay_PIPETX6COMPLIANCE),
    .PIPETX6DATA (delay_PIPETX6DATA),
    .PIPETX6DATAVALID (delay_PIPETX6DATAVALID),
    .PIPETX6ELECIDLE (delay_PIPETX6ELECIDLE),
    .PIPETX6EQCONTROL (delay_PIPETX6EQCONTROL),
    .PIPETX6EQDEEMPH (delay_PIPETX6EQDEEMPH),
    .PIPETX6EQPRESET (delay_PIPETX6EQPRESET),
    .PIPETX6POWERDOWN (delay_PIPETX6POWERDOWN),
    .PIPETX6STARTBLOCK (delay_PIPETX6STARTBLOCK),
    .PIPETX6SYNCHEADER (delay_PIPETX6SYNCHEADER),
    .PIPETX7CHARISK (delay_PIPETX7CHARISK),
    .PIPETX7COMPLIANCE (delay_PIPETX7COMPLIANCE),
    .PIPETX7DATA (delay_PIPETX7DATA),
    .PIPETX7DATAVALID (delay_PIPETX7DATAVALID),
    .PIPETX7ELECIDLE (delay_PIPETX7ELECIDLE),
    .PIPETX7EQCONTROL (delay_PIPETX7EQCONTROL),
    .PIPETX7EQDEEMPH (delay_PIPETX7EQDEEMPH),
    .PIPETX7EQPRESET (delay_PIPETX7EQPRESET),
    .PIPETX7POWERDOWN (delay_PIPETX7POWERDOWN),
    .PIPETX7STARTBLOCK (delay_PIPETX7STARTBLOCK),
    .PIPETX7SYNCHEADER (delay_PIPETX7SYNCHEADER),
    .PIPETXDEEMPH (delay_PIPETXDEEMPH),
    .PIPETXMARGIN (delay_PIPETXMARGIN),
    .PIPETXRATE (delay_PIPETXRATE),
    .PIPETXRCVRDET (delay_PIPETXRCVRDET),
    .PIPETXRESET (delay_PIPETXRESET),
    .PIPETXSWING (delay_PIPETXSWING),
    .PLEQINPROGRESS (delay_PLEQINPROGRESS),
    .PLEQPHASE (delay_PLEQPHASE),
    .PLGEN3PCSRXSLIDE (delay_PLGEN3PCSRXSLIDE),
    .SAXISCCTREADY (delay_SAXISCCTREADY),
    .SAXISRQTREADY (delay_SAXISRQTREADY),
    .CFGCONFIGSPACEENABLE (delay_CFGCONFIGSPACEENABLE),
    .CFGDEVID (delay_CFGDEVID),
    .CFGDSBUSNUMBER (delay_CFGDSBUSNUMBER),
    .CFGDSDEVICENUMBER (delay_CFGDSDEVICENUMBER),
    .CFGDSFUNCTIONNUMBER (delay_CFGDSFUNCTIONNUMBER),
    .CFGDSN (delay_CFGDSN),
    .CFGDSPORTNUMBER (delay_CFGDSPORTNUMBER),
    .CFGERRCORIN (delay_CFGERRCORIN),
    .CFGERRUNCORIN (delay_CFGERRUNCORIN),
    .CFGEXTREADDATA (delay_CFGEXTREADDATA),
    .CFGEXTREADDATAVALID (delay_CFGEXTREADDATAVALID),
    .CFGFCSEL (delay_CFGFCSEL),
    .CFGFLRDONE (delay_CFGFLRDONE),
    .CFGHOTRESETIN (delay_CFGHOTRESETIN),
    .CFGINPUTUPDATEREQUEST (delay_CFGINPUTUPDATEREQUEST),
    .CFGINTERRUPTINT (delay_CFGINTERRUPTINT),
    .CFGINTERRUPTMSIATTR (delay_CFGINTERRUPTMSIATTR),
    .CFGINTERRUPTMSIFUNCTIONNUMBER (delay_CFGINTERRUPTMSIFUNCTIONNUMBER),
    .CFGINTERRUPTMSIINT (delay_CFGINTERRUPTMSIINT),
    .CFGINTERRUPTMSIPENDINGSTATUS (delay_CFGINTERRUPTMSIPENDINGSTATUS),
    .CFGINTERRUPTMSISELECT (delay_CFGINTERRUPTMSISELECT),
    .CFGINTERRUPTMSITPHPRESENT (delay_CFGINTERRUPTMSITPHPRESENT),
    .CFGINTERRUPTMSITPHSTTAG (delay_CFGINTERRUPTMSITPHSTTAG),
    .CFGINTERRUPTMSITPHTYPE (delay_CFGINTERRUPTMSITPHTYPE),
    .CFGINTERRUPTMSIXADDRESS (delay_CFGINTERRUPTMSIXADDRESS),
    .CFGINTERRUPTMSIXDATA (delay_CFGINTERRUPTMSIXDATA),
    .CFGINTERRUPTMSIXINT (delay_CFGINTERRUPTMSIXINT),
    .CFGINTERRUPTPENDING (delay_CFGINTERRUPTPENDING),
    .CFGLINKTRAININGENABLE (delay_CFGLINKTRAININGENABLE),
    .CFGMCUPDATEREQUEST (delay_CFGMCUPDATEREQUEST),
    .CFGMGMTADDR (delay_CFGMGMTADDR),
    .CFGMGMTBYTEENABLE (delay_CFGMGMTBYTEENABLE),
    .CFGMGMTREAD (delay_CFGMGMTREAD),
    .CFGMGMTTYPE1CFGREGACCESS (delay_CFGMGMTTYPE1CFGREGACCESS),
    .CFGMGMTWRITE (delay_CFGMGMTWRITE),
    .CFGMGMTWRITEDATA (delay_CFGMGMTWRITEDATA),
    .CFGMSGTRANSMIT (delay_CFGMSGTRANSMIT),
    .CFGMSGTRANSMITDATA (delay_CFGMSGTRANSMITDATA),
    .CFGMSGTRANSMITTYPE (delay_CFGMSGTRANSMITTYPE),
    .CFGPERFUNCSTATUSCONTROL (delay_CFGPERFUNCSTATUSCONTROL),
    .CFGPERFUNCTIONNUMBER (delay_CFGPERFUNCTIONNUMBER),
    .CFGPERFUNCTIONOUTPUTREQUEST (delay_CFGPERFUNCTIONOUTPUTREQUEST),
    .CFGPOWERSTATECHANGEACK (delay_CFGPOWERSTATECHANGEACK),
    .CFGREQPMTRANSITIONL23READY (delay_CFGREQPMTRANSITIONL23READY),
    .CFGREVID (delay_CFGREVID),
    .CFGSUBSYSID (delay_CFGSUBSYSID),
    .CFGSUBSYSVENDID (delay_CFGSUBSYSVENDID),
    .CFGTPHSTTREADDATA (delay_CFGTPHSTTREADDATA),
    .CFGTPHSTTREADDATAVALID (delay_CFGTPHSTTREADDATAVALID),
    .CFGVENDID (delay_CFGVENDID),
    .CFGVFFLRDONE (delay_CFGVFFLRDONE),
    .CORECLK (delay_CORECLK),
    .CORECLKMICOMPLETIONRAML (delay_CORECLKMICOMPLETIONRAML),
    .CORECLKMICOMPLETIONRAMU (delay_CORECLKMICOMPLETIONRAMU),
    .CORECLKMIREPLAYRAM (delay_CORECLKMIREPLAYRAM),
    .CORECLKMIREQUESTRAM (delay_CORECLKMIREQUESTRAM),
    .DRPADDR (delay_DRPADDR),
    .DRPCLK (delay_DRPCLK),
    .DRPDI (delay_DRPDI),
    .DRPEN (delay_DRPEN),
    .DRPWE (delay_DRPWE),
    .MAXISCQTREADY (delay_MAXISCQTREADY),
    .MAXISRCTREADY (delay_MAXISRCTREADY),
    .MGMTRESETN (delay_MGMTRESETN),
    .MGMTSTICKYRESETN (delay_MGMTSTICKYRESETN),
    .MICOMPLETIONRAMREADDATA (delay_MICOMPLETIONRAMREADDATA),
    .MIREPLAYRAMREADDATA (delay_MIREPLAYRAMREADDATA),
    .MIREQUESTRAMREADDATA (delay_MIREQUESTRAMREADDATA),
    .PCIECQNPREQ (delay_PCIECQNPREQ),
    .PIPECLK (delay_PIPECLK),
    .PIPEEQFS (delay_PIPEEQFS),
    .PIPEEQLF (delay_PIPEEQLF),
    .PIPERESETN (delay_PIPERESETN),
    .PIPERX0CHARISK (delay_PIPERX0CHARISK),
    .PIPERX0DATA (delay_PIPERX0DATA),
    .PIPERX0DATAVALID (delay_PIPERX0DATAVALID),
    .PIPERX0ELECIDLE (delay_PIPERX0ELECIDLE),
    .PIPERX0EQDONE (delay_PIPERX0EQDONE),
    .PIPERX0EQLPADAPTDONE (delay_PIPERX0EQLPADAPTDONE),
    .PIPERX0EQLPLFFSSEL (delay_PIPERX0EQLPLFFSSEL),
    .PIPERX0EQLPNEWTXCOEFFORPRESET (delay_PIPERX0EQLPNEWTXCOEFFORPRESET),
    .PIPERX0PHYSTATUS (delay_PIPERX0PHYSTATUS),
    .PIPERX0STARTBLOCK (delay_PIPERX0STARTBLOCK),
    .PIPERX0STATUS (delay_PIPERX0STATUS),
    .PIPERX0SYNCHEADER (delay_PIPERX0SYNCHEADER),
    .PIPERX0VALID (delay_PIPERX0VALID),
    .PIPERX1CHARISK (delay_PIPERX1CHARISK),
    .PIPERX1DATA (delay_PIPERX1DATA),
    .PIPERX1DATAVALID (delay_PIPERX1DATAVALID),
    .PIPERX1ELECIDLE (delay_PIPERX1ELECIDLE),
    .PIPERX1EQDONE (delay_PIPERX1EQDONE),
    .PIPERX1EQLPADAPTDONE (delay_PIPERX1EQLPADAPTDONE),
    .PIPERX1EQLPLFFSSEL (delay_PIPERX1EQLPLFFSSEL),
    .PIPERX1EQLPNEWTXCOEFFORPRESET (delay_PIPERX1EQLPNEWTXCOEFFORPRESET),
    .PIPERX1PHYSTATUS (delay_PIPERX1PHYSTATUS),
    .PIPERX1STARTBLOCK (delay_PIPERX1STARTBLOCK),
    .PIPERX1STATUS (delay_PIPERX1STATUS),
    .PIPERX1SYNCHEADER (delay_PIPERX1SYNCHEADER),
    .PIPERX1VALID (delay_PIPERX1VALID),
    .PIPERX2CHARISK (delay_PIPERX2CHARISK),
    .PIPERX2DATA (delay_PIPERX2DATA),
    .PIPERX2DATAVALID (delay_PIPERX2DATAVALID),
    .PIPERX2ELECIDLE (delay_PIPERX2ELECIDLE),
    .PIPERX2EQDONE (delay_PIPERX2EQDONE),
    .PIPERX2EQLPADAPTDONE (delay_PIPERX2EQLPADAPTDONE),
    .PIPERX2EQLPLFFSSEL (delay_PIPERX2EQLPLFFSSEL),
    .PIPERX2EQLPNEWTXCOEFFORPRESET (delay_PIPERX2EQLPNEWTXCOEFFORPRESET),
    .PIPERX2PHYSTATUS (delay_PIPERX2PHYSTATUS),
    .PIPERX2STARTBLOCK (delay_PIPERX2STARTBLOCK),
    .PIPERX2STATUS (delay_PIPERX2STATUS),
    .PIPERX2SYNCHEADER (delay_PIPERX2SYNCHEADER),
    .PIPERX2VALID (delay_PIPERX2VALID),
    .PIPERX3CHARISK (delay_PIPERX3CHARISK),
    .PIPERX3DATA (delay_PIPERX3DATA),
    .PIPERX3DATAVALID (delay_PIPERX3DATAVALID),
    .PIPERX3ELECIDLE (delay_PIPERX3ELECIDLE),
    .PIPERX3EQDONE (delay_PIPERX3EQDONE),
    .PIPERX3EQLPADAPTDONE (delay_PIPERX3EQLPADAPTDONE),
    .PIPERX3EQLPLFFSSEL (delay_PIPERX3EQLPLFFSSEL),
    .PIPERX3EQLPNEWTXCOEFFORPRESET (delay_PIPERX3EQLPNEWTXCOEFFORPRESET),
    .PIPERX3PHYSTATUS (delay_PIPERX3PHYSTATUS),
    .PIPERX3STARTBLOCK (delay_PIPERX3STARTBLOCK),
    .PIPERX3STATUS (delay_PIPERX3STATUS),
    .PIPERX3SYNCHEADER (delay_PIPERX3SYNCHEADER),
    .PIPERX3VALID (delay_PIPERX3VALID),
    .PIPERX4CHARISK (delay_PIPERX4CHARISK),
    .PIPERX4DATA (delay_PIPERX4DATA),
    .PIPERX4DATAVALID (delay_PIPERX4DATAVALID),
    .PIPERX4ELECIDLE (delay_PIPERX4ELECIDLE),
    .PIPERX4EQDONE (delay_PIPERX4EQDONE),
    .PIPERX4EQLPADAPTDONE (delay_PIPERX4EQLPADAPTDONE),
    .PIPERX4EQLPLFFSSEL (delay_PIPERX4EQLPLFFSSEL),
    .PIPERX4EQLPNEWTXCOEFFORPRESET (delay_PIPERX4EQLPNEWTXCOEFFORPRESET),
    .PIPERX4PHYSTATUS (delay_PIPERX4PHYSTATUS),
    .PIPERX4STARTBLOCK (delay_PIPERX4STARTBLOCK),
    .PIPERX4STATUS (delay_PIPERX4STATUS),
    .PIPERX4SYNCHEADER (delay_PIPERX4SYNCHEADER),
    .PIPERX4VALID (delay_PIPERX4VALID),
    .PIPERX5CHARISK (delay_PIPERX5CHARISK),
    .PIPERX5DATA (delay_PIPERX5DATA),
    .PIPERX5DATAVALID (delay_PIPERX5DATAVALID),
    .PIPERX5ELECIDLE (delay_PIPERX5ELECIDLE),
    .PIPERX5EQDONE (delay_PIPERX5EQDONE),
    .PIPERX5EQLPADAPTDONE (delay_PIPERX5EQLPADAPTDONE),
    .PIPERX5EQLPLFFSSEL (delay_PIPERX5EQLPLFFSSEL),
    .PIPERX5EQLPNEWTXCOEFFORPRESET (delay_PIPERX5EQLPNEWTXCOEFFORPRESET),
    .PIPERX5PHYSTATUS (delay_PIPERX5PHYSTATUS),
    .PIPERX5STARTBLOCK (delay_PIPERX5STARTBLOCK),
    .PIPERX5STATUS (delay_PIPERX5STATUS),
    .PIPERX5SYNCHEADER (delay_PIPERX5SYNCHEADER),
    .PIPERX5VALID (delay_PIPERX5VALID),
    .PIPERX6CHARISK (delay_PIPERX6CHARISK),
    .PIPERX6DATA (delay_PIPERX6DATA),
    .PIPERX6DATAVALID (delay_PIPERX6DATAVALID),
    .PIPERX6ELECIDLE (delay_PIPERX6ELECIDLE),
    .PIPERX6EQDONE (delay_PIPERX6EQDONE),
    .PIPERX6EQLPADAPTDONE (delay_PIPERX6EQLPADAPTDONE),
    .PIPERX6EQLPLFFSSEL (delay_PIPERX6EQLPLFFSSEL),
    .PIPERX6EQLPNEWTXCOEFFORPRESET (delay_PIPERX6EQLPNEWTXCOEFFORPRESET),
    .PIPERX6PHYSTATUS (delay_PIPERX6PHYSTATUS),
    .PIPERX6STARTBLOCK (delay_PIPERX6STARTBLOCK),
    .PIPERX6STATUS (delay_PIPERX6STATUS),
    .PIPERX6SYNCHEADER (delay_PIPERX6SYNCHEADER),
    .PIPERX6VALID (delay_PIPERX6VALID),
    .PIPERX7CHARISK (delay_PIPERX7CHARISK),
    .PIPERX7DATA (delay_PIPERX7DATA),
    .PIPERX7DATAVALID (delay_PIPERX7DATAVALID),
    .PIPERX7ELECIDLE (delay_PIPERX7ELECIDLE),
    .PIPERX7EQDONE (delay_PIPERX7EQDONE),
    .PIPERX7EQLPADAPTDONE (delay_PIPERX7EQLPADAPTDONE),
    .PIPERX7EQLPLFFSSEL (delay_PIPERX7EQLPLFFSSEL),
    .PIPERX7EQLPNEWTXCOEFFORPRESET (delay_PIPERX7EQLPNEWTXCOEFFORPRESET),
    .PIPERX7PHYSTATUS (delay_PIPERX7PHYSTATUS),
    .PIPERX7STARTBLOCK (delay_PIPERX7STARTBLOCK),
    .PIPERX7STATUS (delay_PIPERX7STATUS),
    .PIPERX7SYNCHEADER (delay_PIPERX7SYNCHEADER),
    .PIPERX7VALID (delay_PIPERX7VALID),
    .PIPETX0EQCOEFF (delay_PIPETX0EQCOEFF),
    .PIPETX0EQDONE (delay_PIPETX0EQDONE),
    .PIPETX1EQCOEFF (delay_PIPETX1EQCOEFF),
    .PIPETX1EQDONE (delay_PIPETX1EQDONE),
    .PIPETX2EQCOEFF (delay_PIPETX2EQCOEFF),
    .PIPETX2EQDONE (delay_PIPETX2EQDONE),
    .PIPETX3EQCOEFF (delay_PIPETX3EQCOEFF),
    .PIPETX3EQDONE (delay_PIPETX3EQDONE),
    .PIPETX4EQCOEFF (delay_PIPETX4EQCOEFF),
    .PIPETX4EQDONE (delay_PIPETX4EQDONE),
    .PIPETX5EQCOEFF (delay_PIPETX5EQCOEFF),
    .PIPETX5EQDONE (delay_PIPETX5EQDONE),
    .PIPETX6EQCOEFF (delay_PIPETX6EQCOEFF),
    .PIPETX6EQDONE (delay_PIPETX6EQDONE),
    .PIPETX7EQCOEFF (delay_PIPETX7EQCOEFF),
    .PIPETX7EQDONE (delay_PIPETX7EQDONE),
    .PLDISABLESCRAMBLER (delay_PLDISABLESCRAMBLER),
    .PLEQRESETEIEOSCOUNT (delay_PLEQRESETEIEOSCOUNT),
    .PLGEN3PCSDISABLE (delay_PLGEN3PCSDISABLE),
    .PLGEN3PCSRXSYNCDONE (delay_PLGEN3PCSRXSYNCDONE),
    .RECCLK (delay_RECCLK),
    .RESETN (delay_RESETN),
    .SAXISCCTDATA (delay_SAXISCCTDATA),
    .SAXISCCTKEEP (delay_SAXISCCTKEEP),
    .SAXISCCTLAST (delay_SAXISCCTLAST),
    .SAXISCCTUSER (delay_SAXISCCTUSER),
    .SAXISCCTVALID (delay_SAXISCCTVALID),
    .SAXISRQTDATA (delay_SAXISRQTDATA),
    .SAXISRQTKEEP (delay_SAXISRQTKEEP),
    .SAXISRQTLAST (delay_SAXISRQTLAST),
    .SAXISRQTUSER (delay_SAXISRQTUSER),
    .SAXISRQTVALID (delay_SAXISRQTVALID),
    .USERCLK (delay_USERCLK)
  );

  specify
    $period (posedge CORECLK, 0:0:0, notifier);
    $period (posedge CORECLKMICOMPLETIONRAML, 0:0:0, notifier);
    $period (posedge CORECLKMICOMPLETIONRAMU, 0:0:0, notifier);
    $period (posedge CORECLKMIREPLAYRAM, 0:0:0, notifier);
    $period (posedge CORECLKMIREQUESTRAM, 0:0:0, notifier);
    $period (posedge DRPCLK, 0:0:0, notifier);
    $period (posedge PIPECLK, 0:0:0, notifier);
    $period (posedge RECCLK, 0:0:0, notifier);
    $period (posedge USERCLK, 0:0:0, notifier);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[0]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[100]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[101]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[102]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[103]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[104]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[105]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[106]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[107]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[108]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[109]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[10]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[110]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[111]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[112]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[113]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[114]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[115]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[116]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[117]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[118]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[119]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[11]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[120]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[121]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[122]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[123]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[124]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[125]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[126]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[127]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[128]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[129]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[12]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[130]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[131]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[132]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[133]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[134]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[135]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[136]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[137]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[138]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[139]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[13]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[140]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[141]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[142]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[143]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[14]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[15]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[16]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[17]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[18]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[19]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[1]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[20]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[21]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[22]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[23]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[24]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[25]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[26]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[27]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[28]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[29]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[2]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[30]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[31]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[32]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[33]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[34]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[35]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[36]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[37]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[38]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[39]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[3]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[40]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[41]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[42]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[43]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[44]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[45]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[46]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[47]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[48]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[49]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[4]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[50]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[51]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[52]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[53]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[54]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[55]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[56]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[57]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[58]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[59]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[5]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[60]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[61]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[62]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[63]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[64]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[65]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[66]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[67]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[68]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[69]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[6]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[70]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[71]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[72]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[73]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[74]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[75]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[76]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[77]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[78]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[79]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[7]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[80]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[81]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[82]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[83]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[84]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[85]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[86]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[87]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[88]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[89]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[8]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[90]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[91]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[92]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[93]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[94]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[95]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[96]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[97]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[98]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[99]);
    $setuphold (posedge CORECLK, negedge MICOMPLETIONRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[9]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[0]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[100]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[101]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[102]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[103]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[104]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[105]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[106]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[107]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[108]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[109]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[10]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[110]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[111]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[112]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[113]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[114]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[115]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[116]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[117]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[118]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[119]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[11]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[120]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[121]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[122]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[123]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[124]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[125]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[126]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[127]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[128]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[129]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[12]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[130]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[131]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[132]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[133]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[134]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[135]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[136]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[137]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[138]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[139]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[13]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[140]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[141]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[142]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[143]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[14]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[15]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[16]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[17]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[18]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[19]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[1]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[20]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[21]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[22]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[23]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[24]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[25]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[26]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[27]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[28]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[29]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[2]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[30]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[31]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[32]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[33]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[34]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[35]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[36]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[37]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[38]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[39]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[3]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[40]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[41]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[42]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[43]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[44]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[45]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[46]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[47]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[48]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[49]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[4]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[50]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[51]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[52]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[53]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[54]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[55]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[56]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[57]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[58]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[59]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[5]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[60]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[61]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[62]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[63]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[64]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[65]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[66]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[67]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[68]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[69]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[6]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[70]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[71]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[72]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[73]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[74]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[75]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[76]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[77]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[78]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[79]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[7]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[80]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[81]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[82]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[83]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[84]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[85]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[86]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[87]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[88]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[89]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[8]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[90]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[91]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[92]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[93]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[94]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[95]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[96]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[97]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[98]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[99]);
    $setuphold (posedge CORECLK, negedge MIREPLAYRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[9]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[0]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[100]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[101]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[102]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[103]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[104]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[105]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[106]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[107]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[108]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[109]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[10]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[110]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[111]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[112]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[113]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[114]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[115]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[116]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[117]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[118]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[119]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[11]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[120]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[121]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[122]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[123]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[124]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[125]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[126]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[127]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[128]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[129]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[12]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[130]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[131]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[132]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[133]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[134]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[135]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[136]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[137]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[138]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[139]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[13]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[140]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[141]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[142]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[143]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[14]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[15]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[16]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[17]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[18]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[19]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[1]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[20]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[21]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[22]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[23]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[24]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[25]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[26]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[27]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[28]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[29]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[2]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[30]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[31]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[32]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[33]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[34]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[35]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[36]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[37]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[38]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[39]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[3]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[40]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[41]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[42]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[43]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[44]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[45]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[46]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[47]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[48]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[49]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[4]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[50]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[51]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[52]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[53]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[54]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[55]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[56]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[57]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[58]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[59]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[5]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[60]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[61]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[62]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[63]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[64]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[65]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[66]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[67]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[68]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[69]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[6]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[70]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[71]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[72]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[73]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[74]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[75]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[76]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[77]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[78]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[79]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[7]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[80]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[81]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[82]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[83]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[84]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[85]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[86]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[87]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[88]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[89]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[8]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[90]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[91]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[92]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[93]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[94]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[95]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[96]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[97]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[98]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[99]);
    $setuphold (posedge CORECLK, negedge MIREQUESTRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[9]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[0]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[100]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[101]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[102]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[103]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[104]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[105]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[106]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[107]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[108]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[109]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[10]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[110]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[111]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[112]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[113]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[114]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[115]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[116]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[117]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[118]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[119]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[11]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[120]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[121]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[122]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[123]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[124]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[125]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[126]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[127]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[128]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[129]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[12]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[130]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[131]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[132]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[133]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[134]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[135]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[136]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[137]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[138]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[139]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[13]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[140]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[141]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[142]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[143]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[14]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[15]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[16]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[17]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[18]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[19]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[1]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[20]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[21]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[22]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[23]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[24]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[25]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[26]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[27]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[28]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[29]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[2]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[30]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[31]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[32]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[33]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[34]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[35]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[36]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[37]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[38]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[39]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[3]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[40]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[41]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[42]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[43]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[44]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[45]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[46]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[47]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[48]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[49]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[4]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[50]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[51]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[52]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[53]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[54]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[55]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[56]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[57]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[58]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[59]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[5]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[60]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[61]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[62]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[63]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[64]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[65]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[66]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[67]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[68]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[69]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[6]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[70]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[71]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[72]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[73]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[74]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[75]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[76]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[77]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[78]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[79]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[7]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[80]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[81]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[82]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[83]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[84]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[85]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[86]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[87]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[88]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[89]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[8]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[90]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[91]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[92]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[93]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[94]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[95]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[96]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[97]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[98]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[99]);
    $setuphold (posedge CORECLK, posedge MICOMPLETIONRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MICOMPLETIONRAMREADDATA[9]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[0]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[100]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[101]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[102]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[103]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[104]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[105]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[106]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[107]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[108]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[109]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[10]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[110]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[111]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[112]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[113]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[114]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[115]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[116]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[117]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[118]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[119]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[11]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[120]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[121]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[122]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[123]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[124]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[125]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[126]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[127]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[128]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[129]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[12]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[130]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[131]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[132]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[133]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[134]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[135]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[136]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[137]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[138]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[139]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[13]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[140]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[141]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[142]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[143]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[14]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[15]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[16]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[17]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[18]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[19]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[1]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[20]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[21]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[22]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[23]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[24]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[25]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[26]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[27]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[28]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[29]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[2]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[30]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[31]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[32]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[33]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[34]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[35]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[36]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[37]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[38]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[39]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[3]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[40]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[41]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[42]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[43]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[44]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[45]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[46]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[47]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[48]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[49]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[4]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[50]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[51]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[52]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[53]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[54]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[55]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[56]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[57]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[58]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[59]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[5]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[60]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[61]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[62]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[63]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[64]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[65]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[66]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[67]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[68]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[69]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[6]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[70]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[71]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[72]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[73]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[74]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[75]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[76]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[77]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[78]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[79]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[7]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[80]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[81]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[82]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[83]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[84]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[85]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[86]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[87]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[88]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[89]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[8]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[90]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[91]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[92]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[93]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[94]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[95]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[96]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[97]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[98]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[99]);
    $setuphold (posedge CORECLK, posedge MIREPLAYRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREPLAYRAMREADDATA[9]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[0]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[100], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[100]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[101], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[101]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[102], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[102]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[103], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[103]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[104], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[104]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[105], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[105]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[106], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[106]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[107], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[107]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[108], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[108]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[109], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[109]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[10]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[110], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[110]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[111], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[111]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[112], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[112]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[113], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[113]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[114], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[114]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[115], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[115]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[116], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[116]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[117], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[117]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[118], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[118]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[119], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[119]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[11]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[120], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[120]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[121], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[121]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[122], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[122]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[123], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[123]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[124], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[124]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[125], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[125]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[126], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[126]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[127], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[127]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[128], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[128]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[129], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[129]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[12]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[130], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[130]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[131], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[131]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[132], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[132]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[133], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[133]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[134], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[134]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[135], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[135]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[136], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[136]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[137], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[137]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[138], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[138]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[139], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[139]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[13]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[140], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[140]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[141], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[141]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[142], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[142]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[143], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[143]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[14]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[15]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[16]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[17]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[18]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[19]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[1]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[20]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[21]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[22]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[23]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[24]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[25]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[26]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[27]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[28]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[29]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[2]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[30]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[31]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[32], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[32]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[33], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[33]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[34], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[34]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[35], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[35]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[36], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[36]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[37], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[37]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[38], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[38]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[39], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[39]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[3]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[40], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[40]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[41], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[41]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[42], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[42]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[43], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[43]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[44], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[44]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[45], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[45]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[46], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[46]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[47], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[47]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[48], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[48]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[49], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[49]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[4]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[50], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[50]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[51], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[51]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[52], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[52]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[53], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[53]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[54], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[54]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[55], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[55]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[56], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[56]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[57], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[57]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[58], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[58]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[59], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[59]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[5]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[60], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[60]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[61], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[61]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[62], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[62]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[63], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[63]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[64], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[64]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[65], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[65]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[66], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[66]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[67], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[67]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[68], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[68]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[69], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[69]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[6]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[70], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[70]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[71], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[71]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[72], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[72]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[73], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[73]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[74], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[74]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[75], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[75]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[76], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[76]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[77], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[77]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[78], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[78]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[79], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[79]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[7]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[80], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[80]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[81], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[81]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[82], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[82]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[83], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[83]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[84], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[84]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[85], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[85]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[86], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[86]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[87], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[87]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[88], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[88]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[89], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[89]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[8]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[90], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[90]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[91], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[91]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[92], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[92]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[93], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[93]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[94], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[94]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[95], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[95]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[96], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[96]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[97], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[97]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[98], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[98]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[99], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[99]);
    $setuphold (posedge CORECLK, posedge MIREQUESTRAMREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_CORECLK, delay_MIREQUESTRAMREADDATA[9]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[0]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[10], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[10]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[1]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[2]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[3]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[4]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[5]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[6]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[7]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[8]);
    $setuphold (posedge DRPCLK, negedge DRPADDR[9], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[9]);
    $setuphold (posedge DRPCLK, negedge DRPDI[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[0]);
    $setuphold (posedge DRPCLK, negedge DRPDI[10], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[10]);
    $setuphold (posedge DRPCLK, negedge DRPDI[11], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[11]);
    $setuphold (posedge DRPCLK, negedge DRPDI[12], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[12]);
    $setuphold (posedge DRPCLK, negedge DRPDI[13], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[13]);
    $setuphold (posedge DRPCLK, negedge DRPDI[14], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[14]);
    $setuphold (posedge DRPCLK, negedge DRPDI[15], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[15]);
    $setuphold (posedge DRPCLK, negedge DRPDI[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[1]);
    $setuphold (posedge DRPCLK, negedge DRPDI[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[2]);
    $setuphold (posedge DRPCLK, negedge DRPDI[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[3]);
    $setuphold (posedge DRPCLK, negedge DRPDI[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[4]);
    $setuphold (posedge DRPCLK, negedge DRPDI[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[5]);
    $setuphold (posedge DRPCLK, negedge DRPDI[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[6]);
    $setuphold (posedge DRPCLK, negedge DRPDI[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[7]);
    $setuphold (posedge DRPCLK, negedge DRPDI[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[8]);
    $setuphold (posedge DRPCLK, negedge DRPDI[9], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[9]);
    $setuphold (posedge DRPCLK, negedge DRPEN, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPEN);
    $setuphold (posedge DRPCLK, negedge DRPWE, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPWE);
    $setuphold (posedge DRPCLK, posedge DRPADDR[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[0]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[10], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[10]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[1]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[2]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[3]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[4]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[5]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[6]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[7]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[8]);
    $setuphold (posedge DRPCLK, posedge DRPADDR[9], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPADDR[9]);
    $setuphold (posedge DRPCLK, posedge DRPDI[0], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[0]);
    $setuphold (posedge DRPCLK, posedge DRPDI[10], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[10]);
    $setuphold (posedge DRPCLK, posedge DRPDI[11], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[11]);
    $setuphold (posedge DRPCLK, posedge DRPDI[12], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[12]);
    $setuphold (posedge DRPCLK, posedge DRPDI[13], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[13]);
    $setuphold (posedge DRPCLK, posedge DRPDI[14], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[14]);
    $setuphold (posedge DRPCLK, posedge DRPDI[15], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[15]);
    $setuphold (posedge DRPCLK, posedge DRPDI[1], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[1]);
    $setuphold (posedge DRPCLK, posedge DRPDI[2], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[2]);
    $setuphold (posedge DRPCLK, posedge DRPDI[3], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[3]);
    $setuphold (posedge DRPCLK, posedge DRPDI[4], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[4]);
    $setuphold (posedge DRPCLK, posedge DRPDI[5], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[5]);
    $setuphold (posedge DRPCLK, posedge DRPDI[6], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[6]);
    $setuphold (posedge DRPCLK, posedge DRPDI[7], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[7]);
    $setuphold (posedge DRPCLK, posedge DRPDI[8], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[8]);
    $setuphold (posedge DRPCLK, posedge DRPDI[9], 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPDI[9]);
    $setuphold (posedge DRPCLK, posedge DRPEN, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPEN);
    $setuphold (posedge DRPCLK, posedge DRPWE, 0:0:0, 0:0:0, notifier,,, delay_DRPCLK, delay_DRPWE);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[0]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[1]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[2]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[3]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[4]);
    $setuphold (posedge PIPECLK, negedge PIPEEQFS[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[5]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[0]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[1]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[2]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[3]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[4]);
    $setuphold (posedge PIPECLK, negedge PIPEEQLF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX0EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX1EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX2EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX3EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX4EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX5EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX6EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, negedge PIPERX7EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX0EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX1EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX2EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX3EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX4EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX5EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX6EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQDONE);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[0]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[10]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[11]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[12]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[13]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[14]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[15]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[16]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[17]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[1]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[2]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[3]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[4]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[5]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[6]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[7]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[8]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[9]);
    $setuphold (posedge PIPECLK, negedge PIPETX7EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQDONE);
    $setuphold (posedge PIPECLK, negedge PLDISABLESCRAMBLER, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDISABLESCRAMBLER);
    $setuphold (posedge PIPECLK, negedge PLEQRESETEIEOSCOUNT, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLEQRESETEIEOSCOUNT);
    $setuphold (posedge PIPECLK, negedge PLGEN3PCSDISABLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLGEN3PCSDISABLE);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[0]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[1]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[2]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[3]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[4]);
    $setuphold (posedge PIPECLK, posedge PIPEEQFS[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQFS[5]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[0]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[1]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[2]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[3]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[4]);
    $setuphold (posedge PIPECLK, posedge PIPEEQLF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPEEQLF[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX0EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX0EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX1EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX1EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX2EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX2EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX3EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX3EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX4EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX4EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX5EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX5EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX6EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX6EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPADAPTDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPADAPTDONE);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPLFFSSEL, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPLFFSSEL);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[0]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[10]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[11]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[12]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[13]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[14]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[15]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[16]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[17]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[1]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[2]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[3]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[4]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[5]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[6]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[7]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[8]);
    $setuphold (posedge PIPECLK, posedge PIPERX7EQLPNEWTXCOEFFORPRESET[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPERX7EQLPNEWTXCOEFFORPRESET[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX0EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX0EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX1EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX1EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX2EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX2EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX3EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX3EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX4EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX4EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX5EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX5EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX6EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX6EQDONE);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[0], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[0]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[10], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[10]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[11], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[11]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[12], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[12]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[13], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[13]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[14], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[14]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[15], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[15]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[16], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[16]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[17], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[17]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[1], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[1]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[2], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[2]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[3], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[3]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[4], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[4]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[5], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[5]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[6], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[6]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[7], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[7]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[8], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[8]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQCOEFF[9], 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQCOEFF[9]);
    $setuphold (posedge PIPECLK, posedge PIPETX7EQDONE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PIPETX7EQDONE);
    $setuphold (posedge PIPECLK, posedge PLDISABLESCRAMBLER, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLDISABLESCRAMBLER);
    $setuphold (posedge PIPECLK, posedge PLEQRESETEIEOSCOUNT, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLEQRESETEIEOSCOUNT);
    $setuphold (posedge PIPECLK, posedge PLGEN3PCSDISABLE, 0:0:0, 0:0:0, notifier,,, delay_PIPECLK, delay_PLGEN3PCSDISABLE);
    $setuphold (posedge RECCLK, negedge PIPERX0CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX0CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX0DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX0ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX0PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX0STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX0STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX0STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX0STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX0SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX0SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX0VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0VALID);
    $setuphold (posedge RECCLK, negedge PIPERX1CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX1CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX1DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX1ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX1PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX1STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX1STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX1STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX1STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX1SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX1SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX1VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1VALID);
    $setuphold (posedge RECCLK, negedge PIPERX2CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX2CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX2DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX2ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX2PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX2STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX2STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX2STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX2STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX2SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX2SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX2VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2VALID);
    $setuphold (posedge RECCLK, negedge PIPERX3CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX3CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX3DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX3ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX3PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX3STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX3STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX3STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX3STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX3SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX3SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX3VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3VALID);
    $setuphold (posedge RECCLK, negedge PIPERX4CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX4CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX4DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX4ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX4PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX4STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX4STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX4STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX4STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX4SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX4SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX4VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4VALID);
    $setuphold (posedge RECCLK, negedge PIPERX5CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX5CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX5DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX5ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX5PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX5STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX5STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX5STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX5STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX5SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX5SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX5VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5VALID);
    $setuphold (posedge RECCLK, negedge PIPERX6CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX6CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX6DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX6ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX6PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX6STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX6STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX6STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX6STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX6SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX6SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX6VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6VALID);
    $setuphold (posedge RECCLK, negedge PIPERX7CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7CHARISK[0]);
    $setuphold (posedge RECCLK, negedge PIPERX7CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7CHARISK[1]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATAVALID);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[0]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[10]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[11]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[12]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[13]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[14]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[15]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[16]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[17]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[18]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[19]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[1]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[20]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[21]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[22]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[23]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[24]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[25]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[26]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[27]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[28]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[29]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[2]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[30]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[31]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[3]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[4]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[5]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[6]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[7]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[8]);
    $setuphold (posedge RECCLK, negedge PIPERX7DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[9]);
    $setuphold (posedge RECCLK, negedge PIPERX7ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7ELECIDLE);
    $setuphold (posedge RECCLK, negedge PIPERX7PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7PHYSTATUS);
    $setuphold (posedge RECCLK, negedge PIPERX7STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STARTBLOCK);
    $setuphold (posedge RECCLK, negedge PIPERX7STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[0]);
    $setuphold (posedge RECCLK, negedge PIPERX7STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[1]);
    $setuphold (posedge RECCLK, negedge PIPERX7STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[2]);
    $setuphold (posedge RECCLK, negedge PIPERX7SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7SYNCHEADER[0]);
    $setuphold (posedge RECCLK, negedge PIPERX7SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7SYNCHEADER[1]);
    $setuphold (posedge RECCLK, negedge PIPERX7VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7VALID);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[0]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[1]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[2]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[3]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[4]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[5]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[6]);
    $setuphold (posedge RECCLK, negedge PLGEN3PCSRXSYNCDONE[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[7]);
    $setuphold (posedge RECCLK, posedge PIPERX0CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX0CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX0DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX0ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX0PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX0STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX0STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX0STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX0STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX0SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX0SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX0VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX0VALID);
    $setuphold (posedge RECCLK, posedge PIPERX1CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX1CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX1DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX1ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX1PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX1STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX1STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX1STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX1STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX1SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX1SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX1VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX1VALID);
    $setuphold (posedge RECCLK, posedge PIPERX2CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX2CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX2DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX2ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX2PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX2STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX2STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX2STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX2STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX2SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX2SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX2VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX2VALID);
    $setuphold (posedge RECCLK, posedge PIPERX3CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX3CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX3DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX3ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX3PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX3STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX3STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX3STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX3STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX3SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX3SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX3VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX3VALID);
    $setuphold (posedge RECCLK, posedge PIPERX4CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX4CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX4DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX4ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX4PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX4STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX4STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX4STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX4STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX4SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX4SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX4VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX4VALID);
    $setuphold (posedge RECCLK, posedge PIPERX5CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX5CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX5DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX5ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX5PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX5STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX5STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX5STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX5STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX5SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX5SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX5VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX5VALID);
    $setuphold (posedge RECCLK, posedge PIPERX6CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX6CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX6DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX6ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX6PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX6STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX6STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX6STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX6STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX6SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX6SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX6VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX6VALID);
    $setuphold (posedge RECCLK, posedge PIPERX7CHARISK[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7CHARISK[0]);
    $setuphold (posedge RECCLK, posedge PIPERX7CHARISK[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7CHARISK[1]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATAVALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATAVALID);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[0]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[10], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[10]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[11], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[11]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[12], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[12]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[13], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[13]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[14], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[14]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[15], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[15]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[16], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[16]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[17], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[17]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[18], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[18]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[19], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[19]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[1]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[20], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[20]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[21], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[21]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[22], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[22]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[23], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[23]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[24], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[24]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[25], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[25]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[26], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[26]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[27], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[27]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[28], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[28]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[29], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[29]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[2]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[30], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[30]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[31], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[31]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[3]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[4]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[5]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[6]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[7]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[8], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[8]);
    $setuphold (posedge RECCLK, posedge PIPERX7DATA[9], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7DATA[9]);
    $setuphold (posedge RECCLK, posedge PIPERX7ELECIDLE, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7ELECIDLE);
    $setuphold (posedge RECCLK, posedge PIPERX7PHYSTATUS, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7PHYSTATUS);
    $setuphold (posedge RECCLK, posedge PIPERX7STARTBLOCK, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STARTBLOCK);
    $setuphold (posedge RECCLK, posedge PIPERX7STATUS[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[0]);
    $setuphold (posedge RECCLK, posedge PIPERX7STATUS[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[1]);
    $setuphold (posedge RECCLK, posedge PIPERX7STATUS[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7STATUS[2]);
    $setuphold (posedge RECCLK, posedge PIPERX7SYNCHEADER[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7SYNCHEADER[0]);
    $setuphold (posedge RECCLK, posedge PIPERX7SYNCHEADER[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7SYNCHEADER[1]);
    $setuphold (posedge RECCLK, posedge PIPERX7VALID, 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PIPERX7VALID);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[0], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[0]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[1], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[1]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[2], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[2]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[3], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[3]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[4], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[4]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[5], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[5]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[6], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[6]);
    $setuphold (posedge RECCLK, posedge PLGEN3PCSRXSYNCDONE[7], 0:0:0, 0:0:0, notifier,,, delay_RECCLK, delay_PLGEN3PCSRXSYNCDONE[7]);
    $setuphold (posedge USERCLK, negedge CFGCONFIGSPACEENABLE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGCONFIGSPACEENABLE);
    $setuphold (posedge USERCLK, negedge CFGDEVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[0]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[10]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[11]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[12]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[13]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[14]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[15]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[1]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[2]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[3]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[4]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[5]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[6]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[7]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[8]);
    $setuphold (posedge USERCLK, negedge CFGDEVID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[9]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[3]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[4]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[5]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[6]);
    $setuphold (posedge USERCLK, negedge CFGDSBUSNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[7]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[3]);
    $setuphold (posedge USERCLK, negedge CFGDSDEVICENUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[4]);
    $setuphold (posedge USERCLK, negedge CFGDSFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGDSFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGDSFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGDSN[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[0]);
    $setuphold (posedge USERCLK, negedge CFGDSN[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[10]);
    $setuphold (posedge USERCLK, negedge CFGDSN[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[11]);
    $setuphold (posedge USERCLK, negedge CFGDSN[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[12]);
    $setuphold (posedge USERCLK, negedge CFGDSN[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[13]);
    $setuphold (posedge USERCLK, negedge CFGDSN[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[14]);
    $setuphold (posedge USERCLK, negedge CFGDSN[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[15]);
    $setuphold (posedge USERCLK, negedge CFGDSN[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[16]);
    $setuphold (posedge USERCLK, negedge CFGDSN[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[17]);
    $setuphold (posedge USERCLK, negedge CFGDSN[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[18]);
    $setuphold (posedge USERCLK, negedge CFGDSN[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[19]);
    $setuphold (posedge USERCLK, negedge CFGDSN[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[1]);
    $setuphold (posedge USERCLK, negedge CFGDSN[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[20]);
    $setuphold (posedge USERCLK, negedge CFGDSN[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[21]);
    $setuphold (posedge USERCLK, negedge CFGDSN[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[22]);
    $setuphold (posedge USERCLK, negedge CFGDSN[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[23]);
    $setuphold (posedge USERCLK, negedge CFGDSN[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[24]);
    $setuphold (posedge USERCLK, negedge CFGDSN[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[25]);
    $setuphold (posedge USERCLK, negedge CFGDSN[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[26]);
    $setuphold (posedge USERCLK, negedge CFGDSN[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[27]);
    $setuphold (posedge USERCLK, negedge CFGDSN[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[28]);
    $setuphold (posedge USERCLK, negedge CFGDSN[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[29]);
    $setuphold (posedge USERCLK, negedge CFGDSN[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[2]);
    $setuphold (posedge USERCLK, negedge CFGDSN[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[30]);
    $setuphold (posedge USERCLK, negedge CFGDSN[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[31]);
    $setuphold (posedge USERCLK, negedge CFGDSN[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[32]);
    $setuphold (posedge USERCLK, negedge CFGDSN[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[33]);
    $setuphold (posedge USERCLK, negedge CFGDSN[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[34]);
    $setuphold (posedge USERCLK, negedge CFGDSN[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[35]);
    $setuphold (posedge USERCLK, negedge CFGDSN[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[36]);
    $setuphold (posedge USERCLK, negedge CFGDSN[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[37]);
    $setuphold (posedge USERCLK, negedge CFGDSN[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[38]);
    $setuphold (posedge USERCLK, negedge CFGDSN[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[39]);
    $setuphold (posedge USERCLK, negedge CFGDSN[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[3]);
    $setuphold (posedge USERCLK, negedge CFGDSN[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[40]);
    $setuphold (posedge USERCLK, negedge CFGDSN[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[41]);
    $setuphold (posedge USERCLK, negedge CFGDSN[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[42]);
    $setuphold (posedge USERCLK, negedge CFGDSN[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[43]);
    $setuphold (posedge USERCLK, negedge CFGDSN[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[44]);
    $setuphold (posedge USERCLK, negedge CFGDSN[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[45]);
    $setuphold (posedge USERCLK, negedge CFGDSN[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[46]);
    $setuphold (posedge USERCLK, negedge CFGDSN[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[47]);
    $setuphold (posedge USERCLK, negedge CFGDSN[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[48]);
    $setuphold (posedge USERCLK, negedge CFGDSN[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[49]);
    $setuphold (posedge USERCLK, negedge CFGDSN[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[4]);
    $setuphold (posedge USERCLK, negedge CFGDSN[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[50]);
    $setuphold (posedge USERCLK, negedge CFGDSN[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[51]);
    $setuphold (posedge USERCLK, negedge CFGDSN[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[52]);
    $setuphold (posedge USERCLK, negedge CFGDSN[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[53]);
    $setuphold (posedge USERCLK, negedge CFGDSN[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[54]);
    $setuphold (posedge USERCLK, negedge CFGDSN[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[55]);
    $setuphold (posedge USERCLK, negedge CFGDSN[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[56]);
    $setuphold (posedge USERCLK, negedge CFGDSN[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[57]);
    $setuphold (posedge USERCLK, negedge CFGDSN[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[58]);
    $setuphold (posedge USERCLK, negedge CFGDSN[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[59]);
    $setuphold (posedge USERCLK, negedge CFGDSN[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[5]);
    $setuphold (posedge USERCLK, negedge CFGDSN[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[60]);
    $setuphold (posedge USERCLK, negedge CFGDSN[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[61]);
    $setuphold (posedge USERCLK, negedge CFGDSN[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[62]);
    $setuphold (posedge USERCLK, negedge CFGDSN[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[63]);
    $setuphold (posedge USERCLK, negedge CFGDSN[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[6]);
    $setuphold (posedge USERCLK, negedge CFGDSN[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[7]);
    $setuphold (posedge USERCLK, negedge CFGDSN[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[8]);
    $setuphold (posedge USERCLK, negedge CFGDSN[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[9]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[3]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[4]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[5]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[6]);
    $setuphold (posedge USERCLK, negedge CFGDSPORTNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[7]);
    $setuphold (posedge USERCLK, negedge CFGERRCORIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGERRCORIN);
    $setuphold (posedge USERCLK, negedge CFGERRUNCORIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGERRUNCORIN);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATAVALID);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[0]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[10]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[11]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[12]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[13]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[14]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[15]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[16]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[17]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[18]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[19]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[1]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[20]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[21]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[22]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[23]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[24]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[25]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[26]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[27]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[28]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[29]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[2]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[30]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[31]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[3]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[4]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[5]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[6]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[7]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[8]);
    $setuphold (posedge USERCLK, negedge CFGEXTREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[9]);
    $setuphold (posedge USERCLK, negedge CFGFCSEL[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[0]);
    $setuphold (posedge USERCLK, negedge CFGFCSEL[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[1]);
    $setuphold (posedge USERCLK, negedge CFGFCSEL[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[2]);
    $setuphold (posedge USERCLK, negedge CFGFLRDONE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFLRDONE[0]);
    $setuphold (posedge USERCLK, negedge CFGFLRDONE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFLRDONE[1]);
    $setuphold (posedge USERCLK, negedge CFGHOTRESETIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGHOTRESETIN);
    $setuphold (posedge USERCLK, negedge CFGINPUTUPDATEREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINPUTUPDATEREQUEST);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTINT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIATTR[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIATTR[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIATTR[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIINT[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[32]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[33]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[34]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[35]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[36]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[37]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[38]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[39]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[40]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[41]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[42]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[43]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[44]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[45]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[46]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[47]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[48]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[49]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[50]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[51]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[52]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[53]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[54]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[55]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[56]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[57]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[58]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[59]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[60]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[61]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[62]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[63]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIPENDINGSTATUS[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSISELECT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHPRESENT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHPRESENT);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHSTTAG[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHTYPE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHTYPE[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSITPHTYPE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHTYPE[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[32]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[33]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[34]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[35]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[36]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[37]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[38]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[39]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[40]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[41]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[42]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[43]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[44]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[45]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[46]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[47]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[48]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[49]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[50]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[51]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[52]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[53]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[54]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[55]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[56]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[57]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[58]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[59]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[60]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[61]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[62]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[63]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXADDRESS[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[10]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[11]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[12]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[13]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[14]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[15]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[16]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[17]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[18]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[19]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[1]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[20]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[21]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[22]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[23]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[24]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[25]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[26]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[27]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[28]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[29]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[2]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[30]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[31]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[3]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[4]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[5]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[6]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[7]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[8]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[9]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTMSIXINT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXINT);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTPENDING[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTPENDING[0]);
    $setuphold (posedge USERCLK, negedge CFGINTERRUPTPENDING[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTPENDING[1]);
    $setuphold (posedge USERCLK, negedge CFGLINKTRAININGENABLE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGLINKTRAININGENABLE);
    $setuphold (posedge USERCLK, negedge CFGMCUPDATEREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMCUPDATEREQUEST);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[0]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[10]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[11]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[12]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[13]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[14]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[15]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[16]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[17]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[18]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[1]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[2]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[3]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[4]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[5]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[6]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[7]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[8]);
    $setuphold (posedge USERCLK, negedge CFGMGMTADDR[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[9]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[0]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[1]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[2]);
    $setuphold (posedge USERCLK, negedge CFGMGMTBYTEENABLE[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[3]);
    $setuphold (posedge USERCLK, negedge CFGMGMTREAD, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTREAD);
    $setuphold (posedge USERCLK, negedge CFGMGMTTYPE1CFGREGACCESS, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTTYPE1CFGREGACCESS);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITE);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[0]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[10]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[11]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[12]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[13]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[14]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[15]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[16]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[17]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[18]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[19]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[1]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[20]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[21]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[22]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[23]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[24]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[25]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[26]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[27]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[28]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[29]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[2]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[30]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[31]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[3]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[4]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[5]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[6]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[7]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[8]);
    $setuphold (posedge USERCLK, negedge CFGMGMTWRITEDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[9]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMIT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMIT);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[0]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[10]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[11]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[12]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[13]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[14]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[15]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[16]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[17]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[18]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[19]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[1]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[20]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[21]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[22]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[23]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[24]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[25]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[26]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[27]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[28]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[29]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[2]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[30]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[31]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[3]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[4]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[5]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[6]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[7]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[8]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[9]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITTYPE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[0]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITTYPE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[1]);
    $setuphold (posedge USERCLK, negedge CFGMSGTRANSMITTYPE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[2]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCSTATUSCONTROL[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[0]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCSTATUSCONTROL[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[1]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCSTATUSCONTROL[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[2]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, negedge CFGPERFUNCTIONOUTPUTREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONOUTPUTREQUEST);
    $setuphold (posedge USERCLK, negedge CFGPOWERSTATECHANGEACK, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPOWERSTATECHANGEACK);
    $setuphold (posedge USERCLK, negedge CFGREQPMTRANSITIONL23READY, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREQPMTRANSITIONL23READY);
    $setuphold (posedge USERCLK, negedge CFGREVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[0]);
    $setuphold (posedge USERCLK, negedge CFGREVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[1]);
    $setuphold (posedge USERCLK, negedge CFGREVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[2]);
    $setuphold (posedge USERCLK, negedge CFGREVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[3]);
    $setuphold (posedge USERCLK, negedge CFGREVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[4]);
    $setuphold (posedge USERCLK, negedge CFGREVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[5]);
    $setuphold (posedge USERCLK, negedge CFGREVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[6]);
    $setuphold (posedge USERCLK, negedge CFGREVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[7]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[0]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[10]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[11]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[12]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[13]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[14]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[15]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[1]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[2]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[3]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[4]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[5]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[6]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[7]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[8]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[9]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[0]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[10]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[11]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[12]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[13]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[14]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[15]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[1]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[2]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[3]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[4]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[5]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[6]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[7]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[8]);
    $setuphold (posedge USERCLK, negedge CFGSUBSYSVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[9]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATAVALID);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[0]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[10]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[11]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[12]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[13]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[14]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[15]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[16]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[17]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[18]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[19]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[1]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[20]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[21]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[22]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[23]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[24]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[25]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[26]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[27]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[28]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[29]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[2]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[30]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[31]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[3]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[4]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[5]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[6]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[7]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[8]);
    $setuphold (posedge USERCLK, negedge CFGTPHSTTREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[9]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[0]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[10]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[11]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[12]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[13]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[14]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[15]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[1]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[2]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[3]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[4]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[5]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[6]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[7]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[8]);
    $setuphold (posedge USERCLK, negedge CFGVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[9]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[0]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[1]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[2]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[3]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[4]);
    $setuphold (posedge USERCLK, negedge CFGVFFLRDONE[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[5]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[0]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[10]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[11]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[12]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[13]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[14]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[15]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[16]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[17]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[18]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[19]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[1]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[20]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[21]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[2]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[3]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[4]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[5]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[6]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[7]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[8]);
    $setuphold (posedge USERCLK, negedge MAXISCQTREADY[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[9]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[0]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[10]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[11]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[12]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[13]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[14]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[15]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[16]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[17]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[18]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[19]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[1]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[20]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[21]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[2]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[3]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[4]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[5]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[6]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[7]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[8]);
    $setuphold (posedge USERCLK, negedge MAXISRCTREADY[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[9]);
    $setuphold (posedge USERCLK, negedge PCIECQNPREQ, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_PCIECQNPREQ);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[0]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[100]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[101]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[102]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[103]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[104]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[105]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[106]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[107]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[108]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[109]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[10]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[110]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[111]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[112]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[113]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[114]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[115]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[116]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[117]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[118]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[119]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[11]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[120]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[121]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[122]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[123]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[124]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[125]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[126]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[127]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[128], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[128]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[129], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[129]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[12]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[130], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[130]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[131], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[131]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[132], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[132]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[133], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[133]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[134], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[134]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[135], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[135]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[136], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[136]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[137], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[137]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[138], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[138]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[139], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[139]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[13]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[140], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[140]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[141], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[141]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[142], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[142]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[143], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[143]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[144], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[144]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[145], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[145]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[146], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[146]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[147], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[147]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[148], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[148]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[149], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[149]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[14]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[150], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[150]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[151], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[151]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[152], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[152]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[153], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[153]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[154], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[154]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[155], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[155]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[156], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[156]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[157], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[157]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[158], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[158]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[159], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[159]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[15]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[160], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[160]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[161], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[161]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[162], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[162]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[163], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[163]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[164], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[164]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[165], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[165]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[166], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[166]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[167], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[167]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[168], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[168]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[169], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[169]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[16]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[170], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[170]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[171], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[171]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[172], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[172]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[173], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[173]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[174], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[174]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[175], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[175]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[176], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[176]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[177], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[177]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[178], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[178]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[179], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[179]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[17]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[180], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[180]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[181], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[181]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[182], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[182]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[183], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[183]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[184], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[184]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[185], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[185]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[186], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[186]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[187], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[187]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[188], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[188]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[189], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[189]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[18]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[190], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[190]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[191], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[191]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[192], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[192]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[193], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[193]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[194], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[194]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[195], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[195]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[196], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[196]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[197], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[197]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[198], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[198]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[199], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[199]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[19]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[1]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[200], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[200]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[201], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[201]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[202], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[202]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[203], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[203]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[204], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[204]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[205], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[205]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[206], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[206]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[207], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[207]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[208], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[208]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[209], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[209]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[20]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[210], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[210]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[211], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[211]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[212], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[212]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[213], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[213]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[214], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[214]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[215], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[215]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[216], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[216]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[217], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[217]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[218], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[218]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[219], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[219]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[21]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[220], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[220]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[221], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[221]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[222], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[222]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[223], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[223]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[224], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[224]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[225], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[225]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[226], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[226]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[227], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[227]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[228], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[228]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[229], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[229]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[22]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[230], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[230]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[231], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[231]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[232], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[232]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[233], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[233]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[234], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[234]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[235], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[235]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[236], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[236]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[237], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[237]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[238], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[238]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[239], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[239]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[23]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[240], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[240]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[241], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[241]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[242], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[242]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[243], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[243]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[244], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[244]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[245], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[245]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[246], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[246]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[247], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[247]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[248], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[248]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[249], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[249]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[24]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[250], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[250]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[251], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[251]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[252], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[252]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[253], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[253]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[254], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[254]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[255], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[255]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[25]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[26]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[27]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[28]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[29]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[2]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[30]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[31]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[32]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[33]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[34]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[35]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[36]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[37]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[38]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[39]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[3]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[40]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[41]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[42]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[43]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[44]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[45]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[46]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[47]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[48]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[49]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[4]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[50]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[51]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[52]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[53]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[54]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[55]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[56]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[57]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[58]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[59]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[5]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[60]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[61]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[62]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[63]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[64]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[65]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[66]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[67]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[68]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[69]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[6]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[70]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[71]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[72]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[73]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[74]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[75]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[76]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[77]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[78]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[79]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[7]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[80]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[81]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[82]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[83]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[84]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[85]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[86]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[87]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[88]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[89]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[8]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[90]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[91]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[92]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[93]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[94]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[95]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[96]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[97]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[98]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[99]);
    $setuphold (posedge USERCLK, negedge SAXISCCTDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[9]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[0]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[1]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[2]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[3]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[4]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[5]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[6]);
    $setuphold (posedge USERCLK, negedge SAXISCCTKEEP[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[7]);
    $setuphold (posedge USERCLK, negedge SAXISCCTLAST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTLAST);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[0]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[10]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[11]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[12]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[13]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[14]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[15]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[16]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[17]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[18]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[19]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[1]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[20]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[21]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[22]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[23]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[24]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[25]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[26]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[27]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[28]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[29]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[2]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[30]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[31]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[32]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[3]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[4]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[5]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[6]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[7]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[8]);
    $setuphold (posedge USERCLK, negedge SAXISCCTUSER[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[9]);
    $setuphold (posedge USERCLK, negedge SAXISCCTVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTVALID);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[0]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[100]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[101]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[102]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[103]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[104]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[105]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[106]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[107]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[108]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[109]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[10]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[110]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[111]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[112]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[113]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[114]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[115]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[116]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[117]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[118]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[119]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[11]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[120]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[121]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[122]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[123]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[124]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[125]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[126]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[127]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[128], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[128]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[129], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[129]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[12]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[130], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[130]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[131], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[131]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[132], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[132]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[133], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[133]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[134], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[134]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[135], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[135]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[136], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[136]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[137], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[137]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[138], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[138]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[139], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[139]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[13]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[140], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[140]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[141], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[141]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[142], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[142]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[143], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[143]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[144], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[144]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[145], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[145]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[146], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[146]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[147], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[147]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[148], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[148]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[149], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[149]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[14]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[150], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[150]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[151], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[151]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[152], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[152]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[153], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[153]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[154], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[154]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[155], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[155]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[156], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[156]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[157], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[157]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[158], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[158]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[159], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[159]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[15]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[160], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[160]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[161], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[161]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[162], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[162]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[163], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[163]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[164], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[164]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[165], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[165]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[166], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[166]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[167], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[167]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[168], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[168]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[169], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[169]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[16]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[170], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[170]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[171], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[171]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[172], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[172]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[173], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[173]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[174], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[174]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[175], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[175]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[176], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[176]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[177], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[177]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[178], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[178]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[179], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[179]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[17]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[180], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[180]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[181], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[181]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[182], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[182]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[183], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[183]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[184], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[184]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[185], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[185]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[186], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[186]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[187], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[187]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[188], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[188]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[189], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[189]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[18]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[190], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[190]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[191], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[191]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[192], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[192]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[193], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[193]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[194], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[194]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[195], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[195]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[196], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[196]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[197], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[197]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[198], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[198]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[199], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[199]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[19]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[1]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[200], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[200]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[201], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[201]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[202], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[202]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[203], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[203]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[204], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[204]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[205], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[205]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[206], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[206]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[207], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[207]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[208], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[208]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[209], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[209]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[20]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[210], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[210]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[211], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[211]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[212], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[212]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[213], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[213]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[214], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[214]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[215], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[215]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[216], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[216]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[217], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[217]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[218], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[218]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[219], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[219]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[21]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[220], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[220]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[221], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[221]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[222], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[222]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[223], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[223]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[224], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[224]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[225], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[225]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[226], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[226]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[227], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[227]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[228], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[228]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[229], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[229]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[22]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[230], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[230]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[231], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[231]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[232], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[232]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[233], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[233]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[234], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[234]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[235], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[235]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[236], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[236]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[237], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[237]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[238], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[238]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[239], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[239]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[23]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[240], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[240]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[241], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[241]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[242], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[242]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[243], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[243]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[244], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[244]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[245], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[245]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[246], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[246]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[247], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[247]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[248], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[248]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[249], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[249]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[24]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[250], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[250]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[251], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[251]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[252], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[252]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[253], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[253]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[254], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[254]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[255], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[255]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[25]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[26]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[27]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[28]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[29]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[2]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[30]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[31]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[32]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[33]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[34]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[35]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[36]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[37]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[38]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[39]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[3]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[40]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[41]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[42]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[43]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[44]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[45]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[46]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[47]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[48]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[49]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[4]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[50]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[51]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[52]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[53]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[54]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[55]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[56]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[57]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[58]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[59]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[5]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[60]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[61]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[62]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[63]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[64]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[65]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[66]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[67]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[68]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[69]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[6]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[70]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[71]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[72]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[73]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[74]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[75]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[76]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[77]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[78]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[79]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[7]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[80]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[81]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[82]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[83]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[84]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[85]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[86]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[87]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[88]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[89]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[8]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[90]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[91]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[92]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[93]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[94]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[95]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[96]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[97]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[98]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[99]);
    $setuphold (posedge USERCLK, negedge SAXISRQTDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[9]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[0]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[1]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[2]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[3]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[4]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[5]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[6]);
    $setuphold (posedge USERCLK, negedge SAXISRQTKEEP[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[7]);
    $setuphold (posedge USERCLK, negedge SAXISRQTLAST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTLAST);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[0]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[10]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[11]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[12]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[13]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[14]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[15]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[16]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[17]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[18]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[19]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[1]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[20]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[21]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[22]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[23]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[24]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[25]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[26]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[27]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[28]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[29]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[2]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[30]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[31]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[32]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[33]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[34]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[35]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[36]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[37]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[38]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[39]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[3]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[40]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[41]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[42]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[43]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[44]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[45]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[46]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[47]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[48]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[49]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[4]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[50]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[51]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[52]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[53]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[54]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[55]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[56]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[57]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[58]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[59]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[5]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[6]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[7]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[8]);
    $setuphold (posedge USERCLK, negedge SAXISRQTUSER[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[9]);
    $setuphold (posedge USERCLK, negedge SAXISRQTVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTVALID);
    $setuphold (posedge USERCLK, posedge CFGCONFIGSPACEENABLE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGCONFIGSPACEENABLE);
    $setuphold (posedge USERCLK, posedge CFGDEVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[0]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[10]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[11]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[12]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[13]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[14]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[15]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[1]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[2]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[3]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[4]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[5]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[6]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[7]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[8]);
    $setuphold (posedge USERCLK, posedge CFGDEVID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDEVID[9]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[3]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[4]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[5]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[6]);
    $setuphold (posedge USERCLK, posedge CFGDSBUSNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSBUSNUMBER[7]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[3]);
    $setuphold (posedge USERCLK, posedge CFGDSDEVICENUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSDEVICENUMBER[4]);
    $setuphold (posedge USERCLK, posedge CFGDSFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGDSFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGDSFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGDSN[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[0]);
    $setuphold (posedge USERCLK, posedge CFGDSN[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[10]);
    $setuphold (posedge USERCLK, posedge CFGDSN[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[11]);
    $setuphold (posedge USERCLK, posedge CFGDSN[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[12]);
    $setuphold (posedge USERCLK, posedge CFGDSN[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[13]);
    $setuphold (posedge USERCLK, posedge CFGDSN[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[14]);
    $setuphold (posedge USERCLK, posedge CFGDSN[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[15]);
    $setuphold (posedge USERCLK, posedge CFGDSN[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[16]);
    $setuphold (posedge USERCLK, posedge CFGDSN[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[17]);
    $setuphold (posedge USERCLK, posedge CFGDSN[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[18]);
    $setuphold (posedge USERCLK, posedge CFGDSN[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[19]);
    $setuphold (posedge USERCLK, posedge CFGDSN[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[1]);
    $setuphold (posedge USERCLK, posedge CFGDSN[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[20]);
    $setuphold (posedge USERCLK, posedge CFGDSN[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[21]);
    $setuphold (posedge USERCLK, posedge CFGDSN[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[22]);
    $setuphold (posedge USERCLK, posedge CFGDSN[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[23]);
    $setuphold (posedge USERCLK, posedge CFGDSN[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[24]);
    $setuphold (posedge USERCLK, posedge CFGDSN[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[25]);
    $setuphold (posedge USERCLK, posedge CFGDSN[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[26]);
    $setuphold (posedge USERCLK, posedge CFGDSN[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[27]);
    $setuphold (posedge USERCLK, posedge CFGDSN[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[28]);
    $setuphold (posedge USERCLK, posedge CFGDSN[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[29]);
    $setuphold (posedge USERCLK, posedge CFGDSN[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[2]);
    $setuphold (posedge USERCLK, posedge CFGDSN[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[30]);
    $setuphold (posedge USERCLK, posedge CFGDSN[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[31]);
    $setuphold (posedge USERCLK, posedge CFGDSN[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[32]);
    $setuphold (posedge USERCLK, posedge CFGDSN[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[33]);
    $setuphold (posedge USERCLK, posedge CFGDSN[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[34]);
    $setuphold (posedge USERCLK, posedge CFGDSN[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[35]);
    $setuphold (posedge USERCLK, posedge CFGDSN[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[36]);
    $setuphold (posedge USERCLK, posedge CFGDSN[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[37]);
    $setuphold (posedge USERCLK, posedge CFGDSN[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[38]);
    $setuphold (posedge USERCLK, posedge CFGDSN[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[39]);
    $setuphold (posedge USERCLK, posedge CFGDSN[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[3]);
    $setuphold (posedge USERCLK, posedge CFGDSN[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[40]);
    $setuphold (posedge USERCLK, posedge CFGDSN[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[41]);
    $setuphold (posedge USERCLK, posedge CFGDSN[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[42]);
    $setuphold (posedge USERCLK, posedge CFGDSN[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[43]);
    $setuphold (posedge USERCLK, posedge CFGDSN[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[44]);
    $setuphold (posedge USERCLK, posedge CFGDSN[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[45]);
    $setuphold (posedge USERCLK, posedge CFGDSN[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[46]);
    $setuphold (posedge USERCLK, posedge CFGDSN[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[47]);
    $setuphold (posedge USERCLK, posedge CFGDSN[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[48]);
    $setuphold (posedge USERCLK, posedge CFGDSN[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[49]);
    $setuphold (posedge USERCLK, posedge CFGDSN[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[4]);
    $setuphold (posedge USERCLK, posedge CFGDSN[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[50]);
    $setuphold (posedge USERCLK, posedge CFGDSN[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[51]);
    $setuphold (posedge USERCLK, posedge CFGDSN[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[52]);
    $setuphold (posedge USERCLK, posedge CFGDSN[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[53]);
    $setuphold (posedge USERCLK, posedge CFGDSN[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[54]);
    $setuphold (posedge USERCLK, posedge CFGDSN[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[55]);
    $setuphold (posedge USERCLK, posedge CFGDSN[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[56]);
    $setuphold (posedge USERCLK, posedge CFGDSN[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[57]);
    $setuphold (posedge USERCLK, posedge CFGDSN[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[58]);
    $setuphold (posedge USERCLK, posedge CFGDSN[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[59]);
    $setuphold (posedge USERCLK, posedge CFGDSN[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[5]);
    $setuphold (posedge USERCLK, posedge CFGDSN[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[60]);
    $setuphold (posedge USERCLK, posedge CFGDSN[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[61]);
    $setuphold (posedge USERCLK, posedge CFGDSN[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[62]);
    $setuphold (posedge USERCLK, posedge CFGDSN[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[63]);
    $setuphold (posedge USERCLK, posedge CFGDSN[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[6]);
    $setuphold (posedge USERCLK, posedge CFGDSN[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[7]);
    $setuphold (posedge USERCLK, posedge CFGDSN[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[8]);
    $setuphold (posedge USERCLK, posedge CFGDSN[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSN[9]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[3]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[4]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[5]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[6]);
    $setuphold (posedge USERCLK, posedge CFGDSPORTNUMBER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGDSPORTNUMBER[7]);
    $setuphold (posedge USERCLK, posedge CFGERRCORIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGERRCORIN);
    $setuphold (posedge USERCLK, posedge CFGERRUNCORIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGERRUNCORIN);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATAVALID);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[0]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[10]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[11]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[12]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[13]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[14]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[15]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[16]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[17]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[18]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[19]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[1]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[20]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[21]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[22]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[23]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[24]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[25]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[26]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[27]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[28]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[29]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[2]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[30]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[31]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[3]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[4]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[5]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[6]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[7]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[8]);
    $setuphold (posedge USERCLK, posedge CFGEXTREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGEXTREADDATA[9]);
    $setuphold (posedge USERCLK, posedge CFGFCSEL[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[0]);
    $setuphold (posedge USERCLK, posedge CFGFCSEL[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[1]);
    $setuphold (posedge USERCLK, posedge CFGFCSEL[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFCSEL[2]);
    $setuphold (posedge USERCLK, posedge CFGFLRDONE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFLRDONE[0]);
    $setuphold (posedge USERCLK, posedge CFGFLRDONE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGFLRDONE[1]);
    $setuphold (posedge USERCLK, posedge CFGHOTRESETIN, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGHOTRESETIN);
    $setuphold (posedge USERCLK, posedge CFGINPUTUPDATEREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINPUTUPDATEREQUEST);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTINT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTINT[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIATTR[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIATTR[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIATTR[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIATTR[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIINT[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIINT[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[32]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[33]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[34]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[35]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[36]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[37]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[38]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[39]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[40]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[41]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[42]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[43]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[44]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[45]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[46]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[47]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[48]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[49]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[50]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[51]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[52]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[53]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[54]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[55]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[56]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[57]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[58]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[59]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[60]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[61]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[62]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[63]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIPENDINGSTATUS[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIPENDINGSTATUS[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSISELECT[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSISELECT[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHPRESENT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHPRESENT);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHSTTAG[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHSTTAG[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHTYPE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHTYPE[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSITPHTYPE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSITPHTYPE[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[32]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[33]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[34]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[35]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[36]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[37]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[38]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[39]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[40]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[41]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[42]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[43]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[44]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[45]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[46]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[47]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[48]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[49]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[50]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[51]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[52]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[53]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[54]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[55]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[56]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[57]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[58]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[59]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[60]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[61]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[62]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[63]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXADDRESS[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXADDRESS[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[10]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[11]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[12]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[13]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[14]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[15]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[16]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[17]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[18]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[19]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[1]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[20]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[21]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[22]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[23]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[24]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[25]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[26]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[27]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[28]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[29]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[2]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[30]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[31]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[3]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[4]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[5]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[6]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[7]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[8]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXDATA[9]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTMSIXINT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTMSIXINT);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTPENDING[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTPENDING[0]);
    $setuphold (posedge USERCLK, posedge CFGINTERRUPTPENDING[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGINTERRUPTPENDING[1]);
    $setuphold (posedge USERCLK, posedge CFGLINKTRAININGENABLE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGLINKTRAININGENABLE);
    $setuphold (posedge USERCLK, posedge CFGMCUPDATEREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMCUPDATEREQUEST);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[0]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[10]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[11]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[12]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[13]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[14]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[15]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[16]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[17]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[18]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[1]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[2]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[3]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[4]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[5]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[6]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[7]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[8]);
    $setuphold (posedge USERCLK, posedge CFGMGMTADDR[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTADDR[9]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[0]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[1]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[2]);
    $setuphold (posedge USERCLK, posedge CFGMGMTBYTEENABLE[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTBYTEENABLE[3]);
    $setuphold (posedge USERCLK, posedge CFGMGMTREAD, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTREAD);
    $setuphold (posedge USERCLK, posedge CFGMGMTTYPE1CFGREGACCESS, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTTYPE1CFGREGACCESS);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITE, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITE);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[0]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[10]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[11]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[12]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[13]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[14]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[15]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[16]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[17]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[18]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[19]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[1]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[20]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[21]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[22]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[23]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[24]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[25]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[26]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[27]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[28]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[29]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[2]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[30]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[31]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[3]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[4]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[5]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[6]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[7]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[8]);
    $setuphold (posedge USERCLK, posedge CFGMGMTWRITEDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMGMTWRITEDATA[9]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMIT, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMIT);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[0]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[10]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[11]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[12]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[13]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[14]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[15]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[16]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[17]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[18]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[19]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[1]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[20]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[21]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[22]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[23]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[24]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[25]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[26]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[27]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[28]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[29]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[2]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[30]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[31]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[3]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[4]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[5]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[6]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[7]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[8]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITDATA[9]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITTYPE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[0]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITTYPE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[1]);
    $setuphold (posedge USERCLK, posedge CFGMSGTRANSMITTYPE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGMSGTRANSMITTYPE[2]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCSTATUSCONTROL[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[0]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCSTATUSCONTROL[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[1]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCSTATUSCONTROL[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCSTATUSCONTROL[2]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONNUMBER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[0]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONNUMBER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[1]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONNUMBER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONNUMBER[2]);
    $setuphold (posedge USERCLK, posedge CFGPERFUNCTIONOUTPUTREQUEST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPERFUNCTIONOUTPUTREQUEST);
    $setuphold (posedge USERCLK, posedge CFGPOWERSTATECHANGEACK, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGPOWERSTATECHANGEACK);
    $setuphold (posedge USERCLK, posedge CFGREQPMTRANSITIONL23READY, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREQPMTRANSITIONL23READY);
    $setuphold (posedge USERCLK, posedge CFGREVID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[0]);
    $setuphold (posedge USERCLK, posedge CFGREVID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[1]);
    $setuphold (posedge USERCLK, posedge CFGREVID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[2]);
    $setuphold (posedge USERCLK, posedge CFGREVID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[3]);
    $setuphold (posedge USERCLK, posedge CFGREVID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[4]);
    $setuphold (posedge USERCLK, posedge CFGREVID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[5]);
    $setuphold (posedge USERCLK, posedge CFGREVID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[6]);
    $setuphold (posedge USERCLK, posedge CFGREVID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGREVID[7]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[0]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[10]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[11]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[12]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[13]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[14]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[15]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[1]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[2]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[3]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[4]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[5]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[6]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[7]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[8]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSID[9]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[0]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[10]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[11]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[12]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[13]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[14]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[15]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[1]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[2]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[3]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[4]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[5]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[6]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[7]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[8]);
    $setuphold (posedge USERCLK, posedge CFGSUBSYSVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGSUBSYSVENDID[9]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATAVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATAVALID);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[0]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[10]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[11]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[12]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[13]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[14]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[15]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[16]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[17]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[18]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[19]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[1]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[20]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[21]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[22]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[23]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[24]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[25]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[26]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[27]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[28]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[29]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[2]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[30]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[31]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[3]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[4]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[5]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[6]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[7]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[8]);
    $setuphold (posedge USERCLK, posedge CFGTPHSTTREADDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGTPHSTTREADDATA[9]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[0]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[10]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[11]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[12]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[13]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[14]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[15]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[1]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[2]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[3]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[4]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[5]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[6]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[7]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[8]);
    $setuphold (posedge USERCLK, posedge CFGVENDID[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVENDID[9]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[0]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[1]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[2]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[3]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[4]);
    $setuphold (posedge USERCLK, posedge CFGVFFLRDONE[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_CFGVFFLRDONE[5]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[0]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[10]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[11]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[12]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[13]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[14]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[15]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[16]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[17]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[18]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[19]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[1]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[20]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[21]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[2]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[3]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[4]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[5]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[6]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[7]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[8]);
    $setuphold (posedge USERCLK, posedge MAXISCQTREADY[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISCQTREADY[9]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[0]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[10]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[11]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[12]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[13]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[14]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[15]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[16]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[17]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[18]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[19]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[1]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[20]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[21]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[2]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[3]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[4]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[5]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[6]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[7]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[8]);
    $setuphold (posedge USERCLK, posedge MAXISRCTREADY[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_MAXISRCTREADY[9]);
    $setuphold (posedge USERCLK, posedge PCIECQNPREQ, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_PCIECQNPREQ);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[0]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[100]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[101]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[102]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[103]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[104]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[105]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[106]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[107]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[108]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[109]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[10]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[110]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[111]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[112]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[113]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[114]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[115]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[116]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[117]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[118]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[119]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[11]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[120]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[121]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[122]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[123]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[124]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[125]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[126]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[127]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[128], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[128]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[129], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[129]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[12]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[130], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[130]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[131], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[131]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[132], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[132]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[133], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[133]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[134], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[134]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[135], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[135]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[136], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[136]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[137], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[137]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[138], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[138]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[139], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[139]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[13]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[140], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[140]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[141], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[141]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[142], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[142]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[143], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[143]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[144], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[144]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[145], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[145]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[146], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[146]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[147], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[147]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[148], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[148]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[149], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[149]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[14]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[150], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[150]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[151], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[151]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[152], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[152]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[153], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[153]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[154], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[154]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[155], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[155]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[156], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[156]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[157], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[157]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[158], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[158]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[159], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[159]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[15]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[160], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[160]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[161], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[161]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[162], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[162]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[163], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[163]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[164], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[164]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[165], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[165]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[166], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[166]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[167], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[167]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[168], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[168]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[169], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[169]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[16]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[170], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[170]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[171], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[171]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[172], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[172]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[173], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[173]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[174], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[174]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[175], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[175]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[176], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[176]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[177], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[177]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[178], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[178]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[179], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[179]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[17]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[180], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[180]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[181], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[181]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[182], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[182]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[183], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[183]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[184], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[184]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[185], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[185]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[186], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[186]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[187], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[187]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[188], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[188]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[189], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[189]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[18]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[190], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[190]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[191], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[191]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[192], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[192]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[193], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[193]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[194], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[194]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[195], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[195]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[196], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[196]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[197], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[197]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[198], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[198]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[199], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[199]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[19]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[1]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[200], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[200]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[201], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[201]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[202], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[202]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[203], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[203]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[204], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[204]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[205], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[205]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[206], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[206]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[207], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[207]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[208], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[208]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[209], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[209]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[20]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[210], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[210]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[211], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[211]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[212], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[212]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[213], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[213]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[214], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[214]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[215], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[215]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[216], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[216]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[217], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[217]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[218], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[218]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[219], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[219]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[21]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[220], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[220]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[221], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[221]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[222], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[222]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[223], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[223]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[224], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[224]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[225], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[225]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[226], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[226]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[227], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[227]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[228], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[228]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[229], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[229]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[22]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[230], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[230]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[231], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[231]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[232], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[232]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[233], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[233]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[234], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[234]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[235], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[235]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[236], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[236]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[237], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[237]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[238], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[238]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[239], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[239]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[23]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[240], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[240]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[241], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[241]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[242], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[242]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[243], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[243]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[244], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[244]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[245], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[245]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[246], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[246]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[247], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[247]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[248], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[248]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[249], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[249]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[24]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[250], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[250]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[251], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[251]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[252], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[252]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[253], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[253]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[254], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[254]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[255], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[255]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[25]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[26]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[27]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[28]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[29]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[2]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[30]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[31]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[32]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[33]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[34]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[35]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[36]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[37]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[38]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[39]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[3]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[40]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[41]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[42]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[43]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[44]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[45]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[46]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[47]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[48]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[49]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[4]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[50]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[51]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[52]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[53]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[54]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[55]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[56]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[57]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[58]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[59]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[5]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[60]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[61]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[62]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[63]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[64]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[65]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[66]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[67]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[68]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[69]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[6]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[70]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[71]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[72]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[73]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[74]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[75]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[76]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[77]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[78]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[79]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[7]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[80]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[81]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[82]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[83]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[84]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[85]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[86]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[87]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[88]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[89]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[8]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[90]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[91]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[92]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[93]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[94]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[95]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[96]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[97]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[98]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[99]);
    $setuphold (posedge USERCLK, posedge SAXISCCTDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTDATA[9]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[0]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[1]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[2]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[3]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[4]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[5]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[6]);
    $setuphold (posedge USERCLK, posedge SAXISCCTKEEP[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTKEEP[7]);
    $setuphold (posedge USERCLK, posedge SAXISCCTLAST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTLAST);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[0]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[10]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[11]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[12]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[13]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[14]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[15]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[16]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[17]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[18]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[19]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[1]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[20]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[21]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[22]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[23]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[24]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[25]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[26]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[27]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[28]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[29]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[2]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[30]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[31]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[32]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[3]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[4]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[5]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[6]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[7]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[8]);
    $setuphold (posedge USERCLK, posedge SAXISCCTUSER[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTUSER[9]);
    $setuphold (posedge USERCLK, posedge SAXISCCTVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISCCTVALID);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[0]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[100], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[100]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[101], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[101]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[102], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[102]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[103], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[103]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[104], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[104]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[105], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[105]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[106], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[106]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[107], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[107]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[108], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[108]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[109], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[109]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[10]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[110], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[110]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[111], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[111]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[112], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[112]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[113], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[113]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[114], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[114]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[115], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[115]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[116], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[116]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[117], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[117]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[118], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[118]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[119], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[119]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[11]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[120], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[120]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[121], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[121]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[122], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[122]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[123], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[123]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[124], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[124]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[125], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[125]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[126], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[126]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[127], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[127]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[128], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[128]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[129], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[129]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[12]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[130], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[130]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[131], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[131]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[132], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[132]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[133], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[133]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[134], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[134]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[135], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[135]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[136], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[136]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[137], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[137]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[138], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[138]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[139], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[139]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[13]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[140], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[140]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[141], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[141]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[142], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[142]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[143], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[143]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[144], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[144]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[145], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[145]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[146], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[146]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[147], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[147]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[148], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[148]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[149], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[149]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[14]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[150], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[150]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[151], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[151]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[152], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[152]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[153], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[153]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[154], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[154]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[155], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[155]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[156], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[156]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[157], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[157]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[158], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[158]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[159], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[159]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[15]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[160], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[160]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[161], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[161]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[162], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[162]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[163], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[163]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[164], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[164]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[165], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[165]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[166], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[166]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[167], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[167]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[168], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[168]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[169], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[169]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[16]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[170], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[170]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[171], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[171]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[172], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[172]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[173], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[173]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[174], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[174]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[175], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[175]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[176], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[176]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[177], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[177]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[178], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[178]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[179], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[179]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[17]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[180], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[180]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[181], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[181]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[182], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[182]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[183], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[183]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[184], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[184]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[185], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[185]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[186], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[186]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[187], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[187]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[188], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[188]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[189], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[189]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[18]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[190], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[190]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[191], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[191]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[192], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[192]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[193], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[193]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[194], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[194]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[195], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[195]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[196], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[196]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[197], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[197]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[198], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[198]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[199], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[199]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[19]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[1]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[200], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[200]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[201], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[201]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[202], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[202]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[203], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[203]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[204], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[204]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[205], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[205]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[206], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[206]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[207], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[207]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[208], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[208]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[209], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[209]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[20]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[210], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[210]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[211], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[211]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[212], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[212]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[213], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[213]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[214], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[214]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[215], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[215]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[216], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[216]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[217], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[217]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[218], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[218]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[219], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[219]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[21]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[220], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[220]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[221], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[221]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[222], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[222]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[223], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[223]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[224], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[224]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[225], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[225]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[226], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[226]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[227], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[227]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[228], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[228]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[229], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[229]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[22]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[230], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[230]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[231], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[231]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[232], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[232]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[233], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[233]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[234], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[234]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[235], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[235]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[236], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[236]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[237], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[237]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[238], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[238]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[239], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[239]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[23]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[240], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[240]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[241], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[241]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[242], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[242]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[243], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[243]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[244], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[244]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[245], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[245]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[246], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[246]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[247], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[247]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[248], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[248]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[249], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[249]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[24]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[250], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[250]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[251], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[251]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[252], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[252]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[253], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[253]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[254], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[254]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[255], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[255]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[25]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[26]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[27]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[28]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[29]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[2]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[30]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[31]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[32]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[33]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[34]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[35]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[36]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[37]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[38]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[39]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[3]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[40]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[41]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[42]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[43]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[44]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[45]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[46]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[47]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[48]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[49]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[4]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[50]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[51]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[52]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[53]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[54]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[55]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[56]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[57]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[58]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[59]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[5]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[60], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[60]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[61], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[61]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[62], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[62]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[63], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[63]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[64], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[64]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[65], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[65]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[66], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[66]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[67], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[67]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[68], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[68]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[69], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[69]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[6]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[70], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[70]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[71], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[71]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[72], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[72]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[73], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[73]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[74], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[74]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[75], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[75]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[76], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[76]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[77], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[77]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[78], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[78]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[79], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[79]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[7]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[80], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[80]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[81], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[81]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[82], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[82]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[83], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[83]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[84], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[84]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[85], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[85]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[86], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[86]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[87], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[87]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[88], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[88]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[89], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[89]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[8]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[90], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[90]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[91], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[91]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[92], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[92]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[93], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[93]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[94], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[94]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[95], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[95]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[96], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[96]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[97], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[97]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[98], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[98]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[99], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[99]);
    $setuphold (posedge USERCLK, posedge SAXISRQTDATA[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTDATA[9]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[0]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[1]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[2]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[3]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[4]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[5]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[6]);
    $setuphold (posedge USERCLK, posedge SAXISRQTKEEP[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTKEEP[7]);
    $setuphold (posedge USERCLK, posedge SAXISRQTLAST, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTLAST);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[0], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[0]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[10], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[10]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[11], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[11]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[12], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[12]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[13], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[13]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[14], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[14]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[15], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[15]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[16], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[16]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[17], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[17]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[18], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[18]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[19], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[19]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[1], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[1]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[20], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[20]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[21], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[21]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[22], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[22]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[23], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[23]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[24], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[24]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[25], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[25]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[26], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[26]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[27], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[27]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[28], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[28]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[29], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[29]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[2], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[2]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[30], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[30]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[31], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[31]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[32], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[32]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[33], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[33]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[34], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[34]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[35], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[35]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[36], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[36]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[37], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[37]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[38], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[38]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[39], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[39]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[3], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[3]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[40], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[40]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[41], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[41]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[42], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[42]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[43], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[43]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[44], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[44]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[45], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[45]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[46], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[46]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[47], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[47]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[48], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[48]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[49], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[49]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[4], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[4]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[50], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[50]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[51], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[51]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[52], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[52]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[53], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[53]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[54], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[54]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[55], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[55]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[56], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[56]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[57], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[57]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[58], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[58]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[59], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[59]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[5], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[5]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[6], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[6]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[7], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[7]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[8], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[8]);
    $setuphold (posedge USERCLK, posedge SAXISRQTUSER[9], 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTUSER[9]);
    $setuphold (posedge USERCLK, posedge SAXISRQTVALID, 0:0:0, 0:0:0, notifier,,, delay_USERCLK, delay_SAXISRQTVALID);
    $width (posedge CORECLK, 0:0:0, 0, notifier);
    $width (posedge CORECLKMICOMPLETIONRAML, 0:0:0, 0, notifier);
    $width (posedge CORECLKMICOMPLETIONRAMU, 0:0:0, 0, notifier);
    $width (posedge CORECLKMIREPLAYRAM, 0:0:0, 0, notifier);
    $width (posedge CORECLKMIREQUESTRAM, 0:0:0, 0, notifier);
    $width (posedge DRPCLK, 0:0:0, 0, notifier);
    $width (posedge PIPECLK, 0:0:0, 0, notifier);
    $width (posedge RECCLK, 0:0:0, 0, notifier);
    $width (posedge USERCLK, 0:0:0, 0, notifier);
    ( CORECLK *> DBGDATAOUT[0]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[10]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[11]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[12]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[13]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[14]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[15]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[1]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[2]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[3]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[4]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[5]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[6]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[7]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[8]) = (100:100:100, 100:100:100);
    ( CORECLK *> DBGDATAOUT[9]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[4]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[5]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[6]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[7]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[8]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSAL[9]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[4]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[5]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[6]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[7]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[8]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADADDRESSBL[9]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADENABLEL[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADENABLEL[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADENABLEL[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMREADENABLEL[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[4]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[5]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[6]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[7]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[8]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSAL[9]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[4]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[5]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[6]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[7]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[8]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEADDRESSBL[9]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[10]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[11]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[12]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[13]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[14]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[15]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[16]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[17]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[18]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[19]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[20]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[21]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[22]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[23]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[24]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[25]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[26]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[27]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[28]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[29]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[30]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[31]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[32]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[33]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[34]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[35]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[36]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[37]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[38]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[39]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[40]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[41]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[42]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[43]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[44]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[45]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[46]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[47]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[48]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[49]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[4]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[50]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[51]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[52]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[53]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[54]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[55]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[56]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[57]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[58]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[59]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[5]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[60]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[61]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[62]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[63]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[64]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[65]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[66]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[67]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[68]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[69]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[6]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[70]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[71]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[7]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[8]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEDATAL[9]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEENABLEL[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEENABLEL[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEENABLEL[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAML *> MICOMPLETIONRAMWRITEENABLEL[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[4]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[5]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[6]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[7]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[8]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSAU[9]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[4]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[5]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[6]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[7]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[8]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADADDRESSBU[9]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADENABLEU[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADENABLEU[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADENABLEU[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMREADENABLEU[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[4]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[5]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[6]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[7]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[8]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSAU[9]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[4]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[5]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[6]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[7]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[8]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEADDRESSBU[9]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[10]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[11]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[12]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[13]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[14]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[15]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[16]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[17]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[18]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[19]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[20]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[21]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[22]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[23]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[24]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[25]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[26]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[27]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[28]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[29]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[30]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[31]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[32]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[33]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[34]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[35]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[36]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[37]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[38]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[39]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[3]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[40]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[41]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[42]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[43]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[44]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[45]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[46]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[47]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[48]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[49]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[4]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[50]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[51]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[52]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[53]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[54]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[55]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[56]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[57]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[58]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[59]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[5]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[60]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[61]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[62]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[63]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[64]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[65]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[66]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[67]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[68]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[69]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[6]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[70]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[71]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[7]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[8]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEDATAU[9]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEENABLEU[0]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEENABLEU[1]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEENABLEU[2]) = (100:100:100, 100:100:100);
    ( CORECLKMICOMPLETIONRAMU *> MICOMPLETIONRAMWRITEENABLEU[3]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[0]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[1]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[2]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[3]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[4]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[5]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[6]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[7]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMADDRESS[8]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMREADENABLE[0]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMREADENABLE[1]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[0]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[100]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[101]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[102]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[103]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[104]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[105]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[106]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[107]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[108]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[109]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[10]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[110]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[111]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[112]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[113]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[114]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[115]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[116]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[117]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[118]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[119]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[11]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[120]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[121]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[122]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[123]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[124]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[125]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[126]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[127]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[128]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[129]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[12]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[130]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[131]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[132]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[133]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[134]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[135]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[136]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[137]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[138]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[139]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[13]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[140]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[141]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[142]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[143]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[14]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[15]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[16]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[17]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[18]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[19]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[1]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[20]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[21]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[22]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[23]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[24]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[25]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[26]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[27]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[28]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[29]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[2]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[30]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[31]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[32]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[33]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[34]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[35]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[36]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[37]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[38]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[39]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[3]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[40]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[41]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[42]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[43]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[44]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[45]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[46]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[47]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[48]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[49]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[4]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[50]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[51]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[52]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[53]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[54]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[55]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[56]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[57]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[58]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[59]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[5]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[60]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[61]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[62]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[63]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[64]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[65]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[66]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[67]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[68]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[69]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[6]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[70]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[71]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[72]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[73]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[74]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[75]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[76]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[77]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[78]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[79]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[7]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[80]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[81]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[82]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[83]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[84]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[85]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[86]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[87]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[88]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[89]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[8]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[90]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[91]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[92]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[93]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[94]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[95]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[96]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[97]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[98]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[99]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEDATA[9]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEENABLE[0]) = (100:100:100, 100:100:100);
    ( CORECLKMIREPLAYRAM *> MIREPLAYRAMWRITEENABLE[1]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[0]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[1]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[2]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[3]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[4]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[5]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[6]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[7]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSA[8]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[0]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[1]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[2]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[3]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[4]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[5]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[6]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[7]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADADDRESSB[8]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADENABLE[0]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADENABLE[1]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADENABLE[2]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMREADENABLE[3]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[0]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[1]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[2]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[3]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[4]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[5]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[6]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[7]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSA[8]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[0]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[1]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[2]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[3]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[4]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[5]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[6]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[7]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEADDRESSB[8]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[0]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[100]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[101]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[102]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[103]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[104]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[105]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[106]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[107]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[108]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[109]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[10]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[110]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[111]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[112]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[113]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[114]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[115]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[116]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[117]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[118]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[119]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[11]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[120]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[121]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[122]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[123]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[124]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[125]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[126]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[127]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[128]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[129]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[12]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[130]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[131]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[132]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[133]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[134]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[135]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[136]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[137]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[138]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[139]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[13]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[140]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[141]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[142]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[143]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[14]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[15]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[16]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[17]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[18]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[19]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[1]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[20]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[21]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[22]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[23]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[24]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[25]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[26]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[27]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[28]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[29]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[2]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[30]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[31]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[32]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[33]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[34]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[35]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[36]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[37]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[38]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[39]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[3]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[40]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[41]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[42]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[43]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[44]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[45]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[46]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[47]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[48]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[49]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[4]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[50]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[51]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[52]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[53]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[54]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[55]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[56]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[57]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[58]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[59]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[5]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[60]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[61]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[62]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[63]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[64]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[65]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[66]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[67]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[68]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[69]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[6]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[70]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[71]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[72]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[73]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[74]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[75]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[76]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[77]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[78]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[79]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[7]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[80]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[81]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[82]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[83]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[84]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[85]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[86]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[87]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[88]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[89]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[8]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[90]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[91]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[92]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[93]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[94]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[95]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[96]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[97]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[98]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[99]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEDATA[9]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEENABLE[0]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEENABLE[1]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEENABLE[2]) = (100:100:100, 100:100:100);
    ( CORECLKMIREQUESTRAM *> MIREQUESTRAMWRITEENABLE[3]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[0]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[10]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[11]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[12]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[13]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[14]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[15]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[1]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[2]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[3]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[4]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[5]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[6]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[7]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[8]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPDO[9]) = (100:100:100, 100:100:100);
    ( DRPCLK *> DRPRDY) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQLPLFFS[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQLPLFFS[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQLPLFFS[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQLPLFFS[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQLPLFFS[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQLPLFFS[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQLPTXPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQLPTXPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQLPTXPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQLPTXPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX0POLARITY) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQLPLFFS[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQLPLFFS[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQLPLFFS[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQLPLFFS[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQLPLFFS[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQLPLFFS[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQLPTXPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQLPTXPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQLPTXPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQLPTXPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX1POLARITY) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQLPLFFS[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQLPLFFS[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQLPLFFS[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQLPLFFS[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQLPLFFS[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQLPLFFS[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQLPTXPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQLPTXPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQLPTXPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQLPTXPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX2POLARITY) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQLPLFFS[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQLPLFFS[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQLPLFFS[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQLPLFFS[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQLPLFFS[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQLPLFFS[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQLPTXPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQLPTXPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQLPTXPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQLPTXPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX3POLARITY) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQLPLFFS[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQLPLFFS[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQLPLFFS[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQLPLFFS[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQLPLFFS[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQLPLFFS[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQLPTXPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQLPTXPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQLPTXPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQLPTXPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX4POLARITY) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQLPLFFS[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQLPLFFS[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQLPLFFS[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQLPLFFS[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQLPLFFS[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQLPLFFS[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQLPTXPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQLPTXPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQLPTXPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQLPTXPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX5POLARITY) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQLPLFFS[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQLPLFFS[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQLPLFFS[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQLPLFFS[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQLPLFFS[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQLPLFFS[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQLPTXPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQLPTXPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQLPTXPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQLPTXPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX6POLARITY) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQLPLFFS[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQLPLFFS[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQLPLFFS[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQLPLFFS[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQLPLFFS[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQLPLFFS[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQLPTXPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQLPTXPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQLPTXPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQLPTXPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPERX7POLARITY) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0CHARISK[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0CHARISK[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0COMPLIANCE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATAVALID) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[10]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[11]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[12]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[13]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[14]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[15]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[16]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[17]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[18]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[19]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[20]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[21]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[22]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[23]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[24]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[25]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[26]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[27]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[28]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[29]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[30]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[31]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[6]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[7]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[8]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0DATA[9]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0ELECIDLE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQDEEMPH[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQDEEMPH[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQDEEMPH[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQDEEMPH[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQDEEMPH[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQDEEMPH[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0EQPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0POWERDOWN[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0POWERDOWN[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0STARTBLOCK) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0SYNCHEADER[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX0SYNCHEADER[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1CHARISK[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1CHARISK[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1COMPLIANCE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATAVALID) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[10]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[11]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[12]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[13]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[14]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[15]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[16]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[17]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[18]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[19]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[20]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[21]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[22]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[23]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[24]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[25]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[26]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[27]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[28]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[29]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[30]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[31]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[6]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[7]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[8]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1DATA[9]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1ELECIDLE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQDEEMPH[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQDEEMPH[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQDEEMPH[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQDEEMPH[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQDEEMPH[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQDEEMPH[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1EQPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1POWERDOWN[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1POWERDOWN[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1STARTBLOCK) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1SYNCHEADER[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX1SYNCHEADER[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2CHARISK[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2CHARISK[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2COMPLIANCE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATAVALID) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[10]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[11]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[12]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[13]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[14]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[15]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[16]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[17]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[18]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[19]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[20]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[21]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[22]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[23]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[24]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[25]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[26]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[27]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[28]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[29]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[30]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[31]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[6]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[7]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[8]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2DATA[9]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2ELECIDLE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQDEEMPH[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQDEEMPH[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQDEEMPH[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQDEEMPH[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQDEEMPH[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQDEEMPH[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2EQPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2POWERDOWN[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2POWERDOWN[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2STARTBLOCK) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2SYNCHEADER[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX2SYNCHEADER[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3CHARISK[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3CHARISK[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3COMPLIANCE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATAVALID) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[10]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[11]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[12]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[13]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[14]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[15]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[16]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[17]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[18]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[19]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[20]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[21]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[22]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[23]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[24]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[25]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[26]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[27]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[28]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[29]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[30]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[31]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[6]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[7]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[8]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3DATA[9]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3ELECIDLE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQDEEMPH[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQDEEMPH[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQDEEMPH[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQDEEMPH[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQDEEMPH[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQDEEMPH[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3EQPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3POWERDOWN[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3POWERDOWN[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3STARTBLOCK) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3SYNCHEADER[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX3SYNCHEADER[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4CHARISK[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4CHARISK[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4COMPLIANCE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATAVALID) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[10]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[11]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[12]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[13]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[14]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[15]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[16]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[17]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[18]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[19]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[20]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[21]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[22]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[23]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[24]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[25]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[26]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[27]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[28]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[29]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[30]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[31]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[6]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[7]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[8]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4DATA[9]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4ELECIDLE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQDEEMPH[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQDEEMPH[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQDEEMPH[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQDEEMPH[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQDEEMPH[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQDEEMPH[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4EQPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4POWERDOWN[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4POWERDOWN[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4STARTBLOCK) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4SYNCHEADER[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX4SYNCHEADER[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5CHARISK[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5CHARISK[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5COMPLIANCE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATAVALID) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[10]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[11]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[12]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[13]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[14]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[15]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[16]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[17]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[18]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[19]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[20]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[21]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[22]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[23]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[24]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[25]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[26]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[27]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[28]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[29]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[30]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[31]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[6]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[7]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[8]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5DATA[9]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5ELECIDLE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQDEEMPH[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQDEEMPH[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQDEEMPH[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQDEEMPH[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQDEEMPH[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQDEEMPH[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5EQPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5POWERDOWN[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5POWERDOWN[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5STARTBLOCK) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5SYNCHEADER[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX5SYNCHEADER[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6CHARISK[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6CHARISK[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6COMPLIANCE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATAVALID) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[10]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[11]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[12]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[13]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[14]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[15]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[16]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[17]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[18]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[19]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[20]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[21]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[22]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[23]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[24]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[25]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[26]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[27]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[28]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[29]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[30]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[31]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[6]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[7]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[8]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6DATA[9]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6ELECIDLE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQDEEMPH[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQDEEMPH[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQDEEMPH[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQDEEMPH[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQDEEMPH[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQDEEMPH[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6EQPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6POWERDOWN[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6POWERDOWN[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6STARTBLOCK) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6SYNCHEADER[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX6SYNCHEADER[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7CHARISK[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7CHARISK[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7COMPLIANCE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATAVALID) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[10]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[11]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[12]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[13]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[14]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[15]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[16]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[17]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[18]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[19]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[20]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[21]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[22]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[23]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[24]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[25]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[26]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[27]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[28]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[29]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[30]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[31]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[6]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[7]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[8]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7DATA[9]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7ELECIDLE) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQCONTROL[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQCONTROL[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQDEEMPH[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQDEEMPH[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQDEEMPH[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQDEEMPH[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQDEEMPH[4]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQDEEMPH[5]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQPRESET[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQPRESET[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQPRESET[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7EQPRESET[3]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7POWERDOWN[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7POWERDOWN[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7STARTBLOCK) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7SYNCHEADER[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETX7SYNCHEADER[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETXDEEMPH) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETXMARGIN[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETXMARGIN[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETXMARGIN[2]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETXRATE[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETXRATE[1]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETXRCVRDET) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETXRESET) = (100:100:100, 100:100:100);
    ( PIPECLK *> PIPETXSWING) = (100:100:100, 100:100:100);
    ( PIPECLK *> PLEQINPROGRESS) = (100:100:100, 100:100:100);
    ( PIPECLK *> PLEQPHASE[0]) = (100:100:100, 100:100:100);
    ( PIPECLK *> PLEQPHASE[1]) = (100:100:100, 100:100:100);
    ( RECCLK *> PLGEN3PCSRXSLIDE[0]) = (100:100:100, 100:100:100);
    ( RECCLK *> PLGEN3PCSRXSLIDE[1]) = (100:100:100, 100:100:100);
    ( RECCLK *> PLGEN3PCSRXSLIDE[2]) = (100:100:100, 100:100:100);
    ( RECCLK *> PLGEN3PCSRXSLIDE[3]) = (100:100:100, 100:100:100);
    ( RECCLK *> PLGEN3PCSRXSLIDE[4]) = (100:100:100, 100:100:100);
    ( RECCLK *> PLGEN3PCSRXSLIDE[5]) = (100:100:100, 100:100:100);
    ( RECCLK *> PLGEN3PCSRXSLIDE[6]) = (100:100:100, 100:100:100);
    ( RECCLK *> PLGEN3PCSRXSLIDE[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGCURRENTSPEED[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGCURRENTSPEED[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGCURRENTSPEED[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGDPASUBSTATECHANGE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGDPASUBSTATECHANGE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGERRCOROUT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGERRFATALOUT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGERRNONFATALOUT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTFUNCTIONNUMBER[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTREADRECEIVED) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTREGISTERNUMBER[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTREGISTERNUMBER[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTREGISTERNUMBER[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTREGISTERNUMBER[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTREGISTERNUMBER[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTREGISTERNUMBER[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTREGISTERNUMBER[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTREGISTERNUMBER[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTREGISTERNUMBER[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTREGISTERNUMBER[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEBYTEENABLE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEBYTEENABLE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEBYTEENABLE[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEBYTEENABLE[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[12]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[13]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[14]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[15]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[16]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[17]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[18]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[19]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[20]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[21]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[22]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[23]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[24]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[25]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[26]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[27]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[28]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[29]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[30]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[31]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITEDATA[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGEXTWRITERECEIVED) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLD[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLH[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLH[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLH[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLH[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLH[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLH[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLH[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCCPLH[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPD[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPH[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPH[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPH[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPH[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPH[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPH[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPH[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCNPH[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPD[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPH[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPH[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPH[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPH[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPH[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPH[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPH[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFCPH[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFLRINPROCESS[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFLRINPROCESS[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONPOWERSTATE[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONSTATUS[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONSTATUS[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONSTATUS[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONSTATUS[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONSTATUS[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONSTATUS[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONSTATUS[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGFUNCTIONSTATUS[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGHOTRESETOUT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINPUTUPDATEDONE) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTAOUTPUT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTBOUTPUT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTCOUTPUT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTDOUTPUT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[12]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[13]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[14]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[15]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[16]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[17]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[18]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[19]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[20]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[21]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[22]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[23]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[24]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[25]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[26]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[27]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[28]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[29]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[30]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[31]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIDATA[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIENABLE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIENABLE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIFAIL) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIMASKUPDATE) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIMMENABLE[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSISENT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIVFENABLE[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXENABLE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXENABLE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXFAIL) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXMASK[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXMASK[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXSENT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFENABLE[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTMSIXVFMASK[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGINTERRUPTSENT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGLINKPOWERSTATE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGLINKPOWERSTATE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGLOCALERROR) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGLTRENABLE) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGLTSSMSTATE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGLTSSMSTATE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGLTSSMSTATE[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGLTSSMSTATE[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGLTSSMSTATE[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGLTSSMSTATE[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMAXPAYLOAD[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMAXPAYLOAD[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMAXPAYLOAD[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMAXREADREQ[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMAXREADREQ[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMAXREADREQ[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMCUPDATEDONE) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[12]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[13]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[14]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[15]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[16]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[17]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[18]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[19]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[20]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[21]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[22]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[23]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[24]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[25]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[26]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[27]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[28]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[29]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[30]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[31]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADDATA[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMGMTREADWRITEDONE) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVED) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDDATA[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDDATA[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDDATA[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDDATA[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDDATA[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDDATA[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDDATA[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDDATA[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDTYPE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDTYPE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDTYPE[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDTYPE[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGRECEIVEDTYPE[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGMSGTRANSMITDONE) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGNEGOTIATEDWIDTH[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGNEGOTIATEDWIDTH[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGNEGOTIATEDWIDTH[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGNEGOTIATEDWIDTH[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGOBFFENABLE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGOBFFENABLE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[12]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[13]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[14]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[15]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCSTATUSDATA[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPERFUNCTIONUPDATEDONE) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPHYLINKDOWN) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPHYLINKSTATUS[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPHYLINKSTATUS[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPLSTATUSCHANGE) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGPOWERSTATECHANGEINTERRUPT) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGRCBSTATUS[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGRCBSTATUS[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHFUNCTIONNUM[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHFUNCTIONNUM[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHFUNCTIONNUM[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHREQUESTERENABLE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHREQUESTERENABLE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTMODE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTMODE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTMODE[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTMODE[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTMODE[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTMODE[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTADDRESS[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTADDRESS[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTADDRESS[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTADDRESS[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTADDRESS[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTREADENABLE) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEBYTEVALID[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEBYTEVALID[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEBYTEVALID[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEBYTEVALID[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[12]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[13]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[14]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[15]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[16]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[17]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[18]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[19]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[20]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[21]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[22]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[23]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[24]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[25]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[26]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[27]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[28]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[29]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[30]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[31]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEDATA[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGTPHSTTWRITEENABLE) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFFLRINPROCESS[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFFLRINPROCESS[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFFLRINPROCESS[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFFLRINPROCESS[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFFLRINPROCESS[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFFLRINPROCESS[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[12]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[13]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[14]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[15]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[16]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[17]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFPOWERSTATE[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFSTATUS[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHREQUESTERENABLE[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[12]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[13]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[14]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[15]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[16]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[17]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> CFGVFTPHSTMODE[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[100]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[101]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[102]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[103]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[104]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[105]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[106]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[107]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[108]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[109]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[110]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[111]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[112]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[113]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[114]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[115]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[116]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[117]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[118]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[119]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[120]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[121]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[122]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[123]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[124]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[125]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[126]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[127]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[128]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[129]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[12]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[130]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[131]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[132]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[133]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[134]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[135]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[136]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[137]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[138]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[139]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[13]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[140]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[141]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[142]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[143]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[144]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[145]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[146]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[147]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[148]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[149]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[14]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[150]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[151]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[152]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[153]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[154]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[155]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[156]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[157]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[158]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[159]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[15]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[160]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[161]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[162]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[163]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[164]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[165]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[166]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[167]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[168]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[169]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[16]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[170]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[171]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[172]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[173]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[174]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[175]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[176]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[177]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[178]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[179]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[17]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[180]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[181]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[182]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[183]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[184]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[185]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[186]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[187]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[188]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[189]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[18]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[190]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[191]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[192]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[193]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[194]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[195]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[196]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[197]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[198]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[199]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[19]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[200]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[201]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[202]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[203]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[204]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[205]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[206]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[207]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[208]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[209]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[20]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[210]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[211]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[212]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[213]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[214]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[215]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[216]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[217]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[218]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[219]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[21]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[220]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[221]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[222]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[223]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[224]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[225]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[226]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[227]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[228]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[229]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[22]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[230]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[231]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[232]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[233]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[234]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[235]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[236]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[237]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[238]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[239]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[23]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[240]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[241]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[242]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[243]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[244]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[245]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[246]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[247]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[248]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[249]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[24]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[250]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[251]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[252]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[253]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[254]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[255]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[25]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[26]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[27]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[28]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[29]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[30]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[31]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[32]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[33]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[34]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[35]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[36]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[37]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[38]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[39]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[40]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[41]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[42]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[43]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[44]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[45]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[46]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[47]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[48]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[49]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[50]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[51]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[52]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[53]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[54]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[55]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[56]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[57]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[58]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[59]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[60]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[61]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[62]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[63]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[64]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[65]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[66]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[67]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[68]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[69]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[70]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[71]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[72]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[73]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[74]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[75]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[76]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[77]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[78]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[79]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[80]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[81]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[82]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[83]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[84]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[85]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[86]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[87]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[88]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[89]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[90]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[91]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[92]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[93]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[94]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[95]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[96]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[97]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[98]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[99]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTDATA[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTKEEP[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTKEEP[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTKEEP[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTKEEP[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTKEEP[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTKEEP[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTKEEP[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTKEEP[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTLAST) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[12]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[13]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[14]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[15]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[16]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[17]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[18]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[19]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[20]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[21]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[22]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[23]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[24]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[25]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[26]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[27]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[28]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[29]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[30]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[31]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[32]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[33]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[34]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[35]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[36]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[37]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[38]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[39]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[40]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[41]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[42]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[43]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[44]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[45]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[46]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[47]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[48]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[49]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[50]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[51]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[52]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[53]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[54]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[55]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[56]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[57]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[58]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[59]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[60]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[61]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[62]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[63]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[64]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[65]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[66]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[67]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[68]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[69]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[70]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[71]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[72]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[73]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[74]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[75]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[76]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[77]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[78]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[79]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[80]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[81]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[82]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[83]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[84]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTUSER[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISCQTVALID) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[100]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[101]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[102]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[103]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[104]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[105]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[106]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[107]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[108]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[109]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[110]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[111]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[112]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[113]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[114]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[115]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[116]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[117]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[118]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[119]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[120]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[121]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[122]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[123]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[124]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[125]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[126]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[127]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[128]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[129]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[12]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[130]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[131]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[132]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[133]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[134]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[135]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[136]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[137]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[138]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[139]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[13]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[140]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[141]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[142]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[143]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[144]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[145]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[146]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[147]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[148]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[149]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[14]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[150]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[151]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[152]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[153]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[154]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[155]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[156]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[157]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[158]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[159]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[15]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[160]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[161]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[162]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[163]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[164]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[165]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[166]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[167]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[168]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[169]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[16]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[170]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[171]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[172]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[173]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[174]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[175]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[176]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[177]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[178]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[179]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[17]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[180]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[181]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[182]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[183]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[184]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[185]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[186]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[187]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[188]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[189]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[18]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[190]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[191]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[192]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[193]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[194]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[195]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[196]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[197]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[198]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[199]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[19]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[200]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[201]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[202]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[203]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[204]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[205]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[206]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[207]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[208]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[209]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[20]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[210]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[211]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[212]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[213]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[214]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[215]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[216]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[217]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[218]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[219]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[21]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[220]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[221]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[222]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[223]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[224]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[225]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[226]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[227]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[228]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[229]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[22]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[230]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[231]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[232]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[233]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[234]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[235]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[236]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[237]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[238]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[239]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[23]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[240]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[241]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[242]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[243]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[244]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[245]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[246]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[247]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[248]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[249]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[24]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[250]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[251]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[252]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[253]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[254]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[255]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[25]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[26]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[27]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[28]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[29]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[30]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[31]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[32]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[33]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[34]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[35]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[36]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[37]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[38]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[39]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[40]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[41]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[42]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[43]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[44]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[45]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[46]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[47]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[48]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[49]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[50]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[51]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[52]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[53]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[54]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[55]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[56]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[57]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[58]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[59]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[60]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[61]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[62]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[63]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[64]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[65]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[66]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[67]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[68]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[69]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[70]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[71]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[72]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[73]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[74]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[75]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[76]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[77]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[78]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[79]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[80]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[81]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[82]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[83]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[84]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[85]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[86]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[87]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[88]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[89]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[90]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[91]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[92]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[93]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[94]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[95]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[96]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[97]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[98]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[99]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTDATA[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTKEEP[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTKEEP[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTKEEP[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTKEEP[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTKEEP[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTKEEP[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTKEEP[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTKEEP[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTLAST) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[10]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[11]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[12]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[13]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[14]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[15]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[16]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[17]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[18]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[19]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[20]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[21]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[22]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[23]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[24]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[25]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[26]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[27]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[28]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[29]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[30]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[31]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[32]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[33]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[34]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[35]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[36]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[37]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[38]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[39]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[40]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[41]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[42]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[43]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[44]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[45]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[46]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[47]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[48]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[49]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[50]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[51]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[52]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[53]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[54]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[55]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[56]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[57]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[58]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[59]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[60]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[61]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[62]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[63]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[64]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[65]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[66]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[67]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[68]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[69]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[6]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[70]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[71]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[72]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[73]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[74]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[7]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[8]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTUSER[9]) = (100:100:100, 100:100:100);
    ( USERCLK *> MAXISRCTVALID) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIECQNPREQCOUNT[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIECQNPREQCOUNT[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIECQNPREQCOUNT[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIECQNPREQCOUNT[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIECQNPREQCOUNT[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIECQNPREQCOUNT[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQSEQNUMVLD) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQSEQNUM[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQSEQNUM[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQSEQNUM[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQSEQNUM[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQTAGAV[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQTAGAV[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQTAGVLD) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQTAG[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQTAG[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQTAG[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQTAG[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQTAG[4]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIERQTAG[5]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIETFCNPDAV[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIETFCNPDAV[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIETFCNPHAV[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> PCIETFCNPHAV[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> SAXISCCTREADY[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> SAXISCCTREADY[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> SAXISCCTREADY[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> SAXISCCTREADY[3]) = (100:100:100, 100:100:100);
    ( USERCLK *> SAXISRQTREADY[0]) = (100:100:100, 100:100:100);
    ( USERCLK *> SAXISRQTREADY[1]) = (100:100:100, 100:100:100);
    ( USERCLK *> SAXISRQTREADY[2]) = (100:100:100, 100:100:100);
    ( USERCLK *> SAXISRQTREADY[3]) = (100:100:100, 100:100:100);

    specparam PATHPULSE$ = 0;
  endspecify
endmodule
