module G_DEPC( q, d, clk, e, p, c );
input c, clk, d, e, p;
output q;
reg q;
parameter initstate = 'b0;

// synthesis translate_off
initial q = initstate;
// synthesis translate_on

always @(posedge clk or posedge p or posedge c)
begin
    if (c == 1'b1)
    begin
        q = 1'b0;
    end
    else if (p == 1'b1)
    begin
        q = 1'b1;
    end
    else if (e == 1'b1)
    begin
        q = d;
    end
end
endmodule

module G_DEC( q, d, clk, e, c );
input c, clk, d, e;
output q;
reg q;
parameter initstate = 'b0;

// synthesis translate_off
initial q = initstate;
// synthesis translate_on

always @(posedge clk or posedge c)
begin
    if (c == 1'b1)
    begin
        q = 1'b0;
    end
    else if (e == 1'b1)
    begin
        q = d;
    end
end
endmodule

module G_DEP( q, d, clk, e, p );
input clk, d, e, p;
output q;
reg q;
parameter initstate = 'b0;

// synthesis translate_off
initial q = initstate;
// synthesis translate_on

always @(posedge clk or posedge p)
begin
     if (p == 1'b1)
     begin
         q = 1'b1;
     end
     else if (e == 1'b1)
     begin
         q = d;
     end
end
endmodule

module G_DE_DEPC( q, d, clk, e, p, c );
input c, clk, d, e, p;
output q;
reg q;
parameter initstate = 'b0;

// synthesis translate_off
initial q = initstate;
// synthesis translate_on

always @(posedge clk or negedge clk or posedge p or posedge c)
begin
    if (c == 1'b1)
    begin
        q = 1'b0;
    end
    else if (p == 1'b1)
    begin
        q = 1'b1;
    end
    else if (e == 1'b1)
    begin
        q = d;
    end
end
endmodule

module G_DE_DEC( q, d, clk, e, c );
input c, clk, d, e;
output q;
reg q;
parameter initstate = 'b0;

// synthesis translate_off
initial q = initstate;
// synthesis translate_on

always @(posedge clk or negedge clk or posedge c)
begin
    if (c == 1'b1)
    begin
        q = 1'b0;
    end
    else if (e == 1'b1)
    begin
        q = d;
    end
end
endmodule

module G_DE_DEP( q, d, clk, e, p );
input clk, d, e, p;
output q;
reg q;
parameter initstate = 'b0;

// synthesis translate_off
initial q = initstate;
// synthesis translate_on

always @(posedge clk or negedge clk or posedge p)
begin
     if (p == 1'b1)
     begin
         q = 1'b1;
     end
     else if (e == 1'b1)
     begin
         q = d;
     end
end
endmodule

module G_TPC ( q, t, clk, p, c );
input clk, p;
output q;
input c, t;
reg q;
parameter initstate = 'b0;

// synthesis translate_off
initial q = initstate;
// synthesis translate_on

always @(posedge clk or posedge p or posedge c)
begin
    if (c == 1'b1)
    begin
        q = 1'b0;
    end
    else if (p == 1'b1)
    begin
        q = 1'b1;
    end
    else if (t == 1'b1)
            q = !q;
end
endmodule

module G_LATPC ( d, p, c, e, q);

  input  d;
  input  p;
  input  c;
  input  e;
  output q;

  wire  d;
  wire  p;
  wire  c;
  wire  e;
  reg   q;
  integer I ;
parameter initstate = 'b0;

// synthesis translate_off
initial q = initstate;
// synthesis translate_on

always @( d or p or c or e) 
begin
    if (c == 1'b1)
        q = 1'b0;
    else if (p == 1'b1)
        q  = 1'b1;
    else if (e == 1'b1)
        q = d;
end
endmodule

module aim_add_sub_2 (ADD_SUB, DATAA0, DATAA1, DATAB0, DATAB1, RESULT0, RESULT1);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAB0;
	input DATAB1;
	output RESULT0;
	output RESULT1;
	wire [1:0] DATAA;
	wire [1:0] DATAB;
	wire [1:0] RESULT;
	assign DATAA = {DATAA1, DATAA0};
	assign DATAB = {DATAB1, DATAB0};
	assign {RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_2 (DATAA0, DATAA1, DATAB0, DATAB1, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAB0;
	input DATAB1;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [1:0] DATAA;
	wire [1:0] DATAB;
	assign DATAA = {DATAA1, DATAA0};
	assign DATAB = {DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_3 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAB0, DATAB1, DATAB2, RESULT0, RESULT1, RESULT2);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	wire [2:0] DATAA;
	wire [2:0] DATAB;
	wire [2:0] RESULT;
	assign DATAA = {DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB2, DATAB1, DATAB0};
	assign {RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_3 (DATAA0, DATAA1, DATAA2, DATAB0, DATAB1, DATAB2, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [2:0] DATAA;
	wire [2:0] DATAB;
	assign DATAA = {DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_4 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAB0, DATAB1, DATAB2, DATAB3, RESULT0, RESULT1, RESULT2, RESULT3);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	wire [3:0] DATAA;
	wire [3:0] DATAB;
	wire [3:0] RESULT;
	assign DATAA = {DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_4 (DATAA0, DATAA1, DATAA2, DATAA3, DATAB0, DATAB1, DATAB2, DATAB3, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [3:0] DATAA;
	wire [3:0] DATAB;
	assign DATAA = {DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_5 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	wire [4:0] DATAA;
	wire [4:0] DATAB;
	wire [4:0] RESULT;
	assign DATAA = {DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_5 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [4:0] DATAA;
	wire [4:0] DATAB;
	assign DATAA = {DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_6 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	wire [5:0] DATAA;
	wire [5:0] DATAB;
	wire [5:0] RESULT;
	assign DATAA = {DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_6 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [5:0] DATAA;
	wire [5:0] DATAB;
	assign DATAA = {DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_7 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	wire [6:0] DATAA;
	wire [6:0] DATAB;
	wire [6:0] RESULT;
	assign DATAA = {DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_7 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [6:0] DATAA;
	wire [6:0] DATAB;
	assign DATAA = {DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_8 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	wire [7:0] DATAA;
	wire [7:0] DATAB;
	wire [7:0] RESULT;
	assign DATAA = {DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_8 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [7:0] DATAA;
	wire [7:0] DATAB;
	assign DATAA = {DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_9 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	wire [8:0] DATAA;
	wire [8:0] DATAB;
	wire [8:0] RESULT;
	assign DATAA = {DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_9 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [8:0] DATAA;
	wire [8:0] DATAB;
	assign DATAA = {DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_10 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	wire [9:0] DATAA;
	wire [9:0] DATAB;
	wire [9:0] RESULT;
	assign DATAA = {DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_10 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [9:0] DATAA;
	wire [9:0] DATAB;
	assign DATAA = {DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_11 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	wire [10:0] DATAA;
	wire [10:0] DATAB;
	wire [10:0] RESULT;
	assign DATAA = {DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_11 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [10:0] DATAA;
	wire [10:0] DATAB;
	assign DATAA = {DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_12 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	wire [11:0] DATAA;
	wire [11:0] DATAB;
	wire [11:0] RESULT;
	assign DATAA = {DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_12 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [11:0] DATAA;
	wire [11:0] DATAB;
	assign DATAA = {DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_13 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	wire [12:0] DATAA;
	wire [12:0] DATAB;
	wire [12:0] RESULT;
	assign DATAA = {DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_13 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [12:0] DATAA;
	wire [12:0] DATAB;
	assign DATAA = {DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_14 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	wire [13:0] DATAA;
	wire [13:0] DATAB;
	wire [13:0] RESULT;
	assign DATAA = {DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_14 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [13:0] DATAA;
	wire [13:0] DATAB;
	assign DATAA = {DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_15 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	wire [14:0] DATAA;
	wire [14:0] DATAB;
	wire [14:0] RESULT;
	assign DATAA = {DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_15 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [14:0] DATAA;
	wire [14:0] DATAB;
	assign DATAA = {DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_16 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	wire [15:0] DATAA;
	wire [15:0] DATAB;
	wire [15:0] RESULT;
	assign DATAA = {DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_16 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [15:0] DATAA;
	wire [15:0] DATAB;
	assign DATAA = {DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_17 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	wire [16:0] DATAA;
	wire [16:0] DATAB;
	wire [16:0] RESULT;
	assign DATAA = {DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_17 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [16:0] DATAA;
	wire [16:0] DATAB;
	assign DATAA = {DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_18 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	wire [17:0] DATAA;
	wire [17:0] DATAB;
	wire [17:0] RESULT;
	assign DATAA = {DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_18 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [17:0] DATAA;
	wire [17:0] DATAB;
	assign DATAA = {DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_19 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	wire [18:0] DATAA;
	wire [18:0] DATAB;
	wire [18:0] RESULT;
	assign DATAA = {DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_19 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [18:0] DATAA;
	wire [18:0] DATAB;
	assign DATAA = {DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_20 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	wire [19:0] DATAA;
	wire [19:0] DATAB;
	wire [19:0] RESULT;
	assign DATAA = {DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_20 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [19:0] DATAA;
	wire [19:0] DATAB;
	assign DATAA = {DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_21 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19, RESULT20);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	output RESULT20;
	wire [20:0] DATAA;
	wire [20:0] DATAB;
	wire [20:0] RESULT;
	assign DATAA = {DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_21 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [20:0] DATAA;
	wire [20:0] DATAB;
	assign DATAA = {DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_22 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19, RESULT20, RESULT21);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	output RESULT20;
	output RESULT21;
	wire [21:0] DATAA;
	wire [21:0] DATAB;
	wire [21:0] RESULT;
	assign DATAA = {DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT21, RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_22 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [21:0] DATAA;
	wire [21:0] DATAB;
	assign DATAA = {DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_23 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19, RESULT20, RESULT21, RESULT22);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	output RESULT20;
	output RESULT21;
	output RESULT22;
	wire [22:0] DATAA;
	wire [22:0] DATAB;
	wire [22:0] RESULT;
	assign DATAA = {DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT22, RESULT21, RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_23 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [22:0] DATAA;
	wire [22:0] DATAB;
	assign DATAA = {DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_24 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19, RESULT20, RESULT21, RESULT22, RESULT23);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	output RESULT20;
	output RESULT21;
	output RESULT22;
	output RESULT23;
	wire [23:0] DATAA;
	wire [23:0] DATAB;
	wire [23:0] RESULT;
	assign DATAA = {DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT23, RESULT22, RESULT21, RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_24 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [23:0] DATAA;
	wire [23:0] DATAB;
	assign DATAA = {DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_25 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19, RESULT20, RESULT21, RESULT22, RESULT23, RESULT24);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	output RESULT20;
	output RESULT21;
	output RESULT22;
	output RESULT23;
	output RESULT24;
	wire [24:0] DATAA;
	wire [24:0] DATAB;
	wire [24:0] RESULT;
	assign DATAA = {DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT24, RESULT23, RESULT22, RESULT21, RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_25 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [24:0] DATAA;
	wire [24:0] DATAB;
	assign DATAA = {DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_26 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19, RESULT20, RESULT21, RESULT22, RESULT23, RESULT24, RESULT25);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	output RESULT20;
	output RESULT21;
	output RESULT22;
	output RESULT23;
	output RESULT24;
	output RESULT25;
	wire [25:0] DATAA;
	wire [25:0] DATAB;
	wire [25:0] RESULT;
	assign DATAA = {DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT25, RESULT24, RESULT23, RESULT22, RESULT21, RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_26 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [25:0] DATAA;
	wire [25:0] DATAB;
	assign DATAA = {DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_27 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAA26, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, DATAB26, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19, RESULT20, RESULT21, RESULT22, RESULT23, RESULT24, RESULT25, RESULT26);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAA26;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	input DATAB26;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	output RESULT20;
	output RESULT21;
	output RESULT22;
	output RESULT23;
	output RESULT24;
	output RESULT25;
	output RESULT26;
	wire [26:0] DATAA;
	wire [26:0] DATAB;
	wire [26:0] RESULT;
	assign DATAA = {DATAA26, DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB26, DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT26, RESULT25, RESULT24, RESULT23, RESULT22, RESULT21, RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_27 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAA26, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, DATAB26, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAA26;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	input DATAB26;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [26:0] DATAA;
	wire [26:0] DATAB;
	assign DATAA = {DATAA26, DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB26, DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_28 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAA26, DATAA27, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, DATAB26, DATAB27, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19, RESULT20, RESULT21, RESULT22, RESULT23, RESULT24, RESULT25, RESULT26, RESULT27);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAA26;
	input DATAA27;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	input DATAB26;
	input DATAB27;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	output RESULT20;
	output RESULT21;
	output RESULT22;
	output RESULT23;
	output RESULT24;
	output RESULT25;
	output RESULT26;
	output RESULT27;
	wire [27:0] DATAA;
	wire [27:0] DATAB;
	wire [27:0] RESULT;
	assign DATAA = {DATAA27, DATAA26, DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB27, DATAB26, DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT27, RESULT26, RESULT25, RESULT24, RESULT23, RESULT22, RESULT21, RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_28 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAA26, DATAA27, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, DATAB26, DATAB27, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAA26;
	input DATAA27;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	input DATAB26;
	input DATAB27;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [27:0] DATAA;
	wire [27:0] DATAB;
	assign DATAA = {DATAA27, DATAA26, DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB27, DATAB26, DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_29 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAA26, DATAA27, DATAA28, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, DATAB26, DATAB27, DATAB28, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19, RESULT20, RESULT21, RESULT22, RESULT23, RESULT24, RESULT25, RESULT26, RESULT27, RESULT28);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAA26;
	input DATAA27;
	input DATAA28;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	input DATAB26;
	input DATAB27;
	input DATAB28;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	output RESULT20;
	output RESULT21;
	output RESULT22;
	output RESULT23;
	output RESULT24;
	output RESULT25;
	output RESULT26;
	output RESULT27;
	output RESULT28;
	wire [28:0] DATAA;
	wire [28:0] DATAB;
	wire [28:0] RESULT;
	assign DATAA = {DATAA28, DATAA27, DATAA26, DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB28, DATAB27, DATAB26, DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT28, RESULT27, RESULT26, RESULT25, RESULT24, RESULT23, RESULT22, RESULT21, RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_29 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAA26, DATAA27, DATAA28, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, DATAB26, DATAB27, DATAB28, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAA26;
	input DATAA27;
	input DATAA28;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	input DATAB26;
	input DATAB27;
	input DATAB28;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [28:0] DATAA;
	wire [28:0] DATAB;
	assign DATAA = {DATAA28, DATAA27, DATAA26, DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB28, DATAB27, DATAB26, DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_30 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAA26, DATAA27, DATAA28, DATAA29, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, DATAB26, DATAB27, DATAB28, DATAB29, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19, RESULT20, RESULT21, RESULT22, RESULT23, RESULT24, RESULT25, RESULT26, RESULT27, RESULT28, RESULT29);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAA26;
	input DATAA27;
	input DATAA28;
	input DATAA29;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	input DATAB26;
	input DATAB27;
	input DATAB28;
	input DATAB29;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	output RESULT20;
	output RESULT21;
	output RESULT22;
	output RESULT23;
	output RESULT24;
	output RESULT25;
	output RESULT26;
	output RESULT27;
	output RESULT28;
	output RESULT29;
	wire [29:0] DATAA;
	wire [29:0] DATAB;
	wire [29:0] RESULT;
	assign DATAA = {DATAA29, DATAA28, DATAA27, DATAA26, DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB29, DATAB28, DATAB27, DATAB26, DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT29, RESULT28, RESULT27, RESULT26, RESULT25, RESULT24, RESULT23, RESULT22, RESULT21, RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_30 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAA26, DATAA27, DATAA28, DATAA29, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, DATAB26, DATAB27, DATAB28, DATAB29, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAA26;
	input DATAA27;
	input DATAA28;
	input DATAA29;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	input DATAB26;
	input DATAB27;
	input DATAB28;
	input DATAB29;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [29:0] DATAA;
	wire [29:0] DATAB;
	assign DATAA = {DATAA29, DATAA28, DATAA27, DATAA26, DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB29, DATAB28, DATAB27, DATAB26, DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

module aim_add_sub_31 (ADD_SUB, DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAA26, DATAA27, DATAA28, DATAA29, DATAA30, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, DATAB26, DATAB27, DATAB28, DATAB29, DATAB30, RESULT0, RESULT1, RESULT2, RESULT3, RESULT4, RESULT5, RESULT6, RESULT7, RESULT8, RESULT9, RESULT10, RESULT11, RESULT12, RESULT13, RESULT14, RESULT15, RESULT16, RESULT17, RESULT18, RESULT19, RESULT20, RESULT21, RESULT22, RESULT23, RESULT24, RESULT25, RESULT26, RESULT27, RESULT28, RESULT29, RESULT30);
	input ADD_SUB;
	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAA26;
	input DATAA27;
	input DATAA28;
	input DATAA29;
	input DATAA30;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	input DATAB26;
	input DATAB27;
	input DATAB28;
	input DATAB29;
	input DATAB30;
	output RESULT0;
	output RESULT1;
	output RESULT2;
	output RESULT3;
	output RESULT4;
	output RESULT5;
	output RESULT6;
	output RESULT7;
	output RESULT8;
	output RESULT9;
	output RESULT10;
	output RESULT11;
	output RESULT12;
	output RESULT13;
	output RESULT14;
	output RESULT15;
	output RESULT16;
	output RESULT17;
	output RESULT18;
	output RESULT19;
	output RESULT20;
	output RESULT21;
	output RESULT22;
	output RESULT23;
	output RESULT24;
	output RESULT25;
	output RESULT26;
	output RESULT27;
	output RESULT28;
	output RESULT29;
	output RESULT30;
	wire [30:0] DATAA;
	wire [30:0] DATAB;
	wire [30:0] RESULT;
	assign DATAA = {DATAA30, DATAA29, DATAA28, DATAA27, DATAA26, DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB30, DATAB29, DATAB28, DATAB27, DATAB26, DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign {RESULT30, RESULT29, RESULT28, RESULT27, RESULT26, RESULT25, RESULT24, RESULT23, RESULT22, RESULT21, RESULT20, RESULT19, RESULT18, RESULT17, RESULT16, RESULT15, RESULT14, RESULT13, RESULT12, RESULT11, RESULT10, RESULT9, RESULT8, RESULT7, RESULT6, RESULT5, RESULT4, RESULT3, RESULT2, RESULT1, RESULT0} = RESULT;
	assign RESULT = (ADD_SUB == 'b1) ? DATAA+DATAB : DATAA-DATAB;
endmodule

module aim_compare_31 (DATAA0, DATAA1, DATAA2, DATAA3, DATAA4, DATAA5, DATAA6, DATAA7, DATAA8, DATAA9, DATAA10, DATAA11, DATAA12, DATAA13, DATAA14, DATAA15, DATAA16, DATAA17, DATAA18, DATAA19, DATAA20, DATAA21, DATAA22, DATAA23, DATAA24, DATAA25, DATAA26, DATAA27, DATAA28, DATAA29, DATAA30, DATAB0, DATAB1, DATAB2, DATAB3, DATAB4, DATAB5, DATAB6, DATAB7, DATAB8, DATAB9, DATAB10, DATAB11, DATAB12, DATAB13, DATAB14, DATAB15, DATAB16, DATAB17, DATAB18, DATAB19, DATAB20, DATAB21, DATAB22, DATAB23, DATAB24, DATAB25, DATAB26, DATAB27, DATAB28, DATAB29, DATAB30, AEB, ANEB, AGB, AGEB, ALB, ALEB);	input DATAA0;
	input DATAA1;
	input DATAA2;
	input DATAA3;
	input DATAA4;
	input DATAA5;
	input DATAA6;
	input DATAA7;
	input DATAA8;
	input DATAA9;
	input DATAA10;
	input DATAA11;
	input DATAA12;
	input DATAA13;
	input DATAA14;
	input DATAA15;
	input DATAA16;
	input DATAA17;
	input DATAA18;
	input DATAA19;
	input DATAA20;
	input DATAA21;
	input DATAA22;
	input DATAA23;
	input DATAA24;
	input DATAA25;
	input DATAA26;
	input DATAA27;
	input DATAA28;
	input DATAA29;
	input DATAA30;
	input DATAB0;
	input DATAB1;
	input DATAB2;
	input DATAB3;
	input DATAB4;
	input DATAB5;
	input DATAB6;
	input DATAB7;
	input DATAB8;
	input DATAB9;
	input DATAB10;
	input DATAB11;
	input DATAB12;
	input DATAB13;
	input DATAB14;
	input DATAB15;
	input DATAB16;
	input DATAB17;
	input DATAB18;
	input DATAB19;
	input DATAB20;
	input DATAB21;
	input DATAB22;
	input DATAB23;
	input DATAB24;
	input DATAB25;
	input DATAB26;
	input DATAB27;
	input DATAB28;
	input DATAB29;
	input DATAB30;
	output AEB, ANEB, AGB, AGEB, ALB, ALEB;
	wire [30:0] DATAA;
	wire [30:0] DATAB;
	assign DATAA = {DATAA30, DATAA29, DATAA28, DATAA27, DATAA26, DATAA25, DATAA24, DATAA23, DATAA22, DATAA21, DATAA20, DATAA19, DATAA18, DATAA17, DATAA16, DATAA15, DATAA14, DATAA13, DATAA12, DATAA11, DATAA10, DATAA9, DATAA8, DATAA7, DATAA6, DATAA5, DATAA4, DATAA3, DATAA2, DATAA1, DATAA0};
	assign DATAB = {DATAB30, DATAB29, DATAB28, DATAB27, DATAB26, DATAB25, DATAB24, DATAB23, DATAB22, DATAB21, DATAB20, DATAB19, DATAB18, DATAB17, DATAB16, DATAB15, DATAB14, DATAB13, DATAB12, DATAB11, DATAB10, DATAB9, DATAB8, DATAB7, DATAB6, DATAB5, DATAB4, DATAB3, DATAB2, DATAB1, DATAB0};
	assign AEB = (DATAA == DATAB) ? 'b1 : 'b0;
	assign ANEB = (DATAA != DATAB) ? 'b1 : 'b0;
	assign AGB = (DATAA > DATAB) ? 'b1 : 'b0;
	assign AGEB = (DATAA >= DATAB) ? 'b1 : 'b0;
	assign ALB = (DATAA < DATAB) ? 'b1 : 'b0;
	assign ALEB = (DATAA <= DATAB) ? 'b1 : 'b0;
endmodule

